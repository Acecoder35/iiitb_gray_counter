magic
tech sky130A
magscale 1 2
timestamp 1670837674
<< viali >>
rect 1777 9129 1811 9163
rect 6745 9129 6779 9163
rect 8033 9129 8067 9163
rect 1593 8925 1627 8959
rect 6561 8925 6595 8959
rect 7849 8925 7883 8959
rect 1777 8585 1811 8619
rect 1593 8449 1627 8483
rect 4445 7837 4479 7871
rect 4905 7837 4939 7871
rect 5089 7837 5123 7871
rect 7849 7837 7883 7871
rect 4261 7701 4295 7735
rect 4997 7701 5031 7735
rect 8033 7701 8067 7735
rect 1593 7497 1627 7531
rect 5549 7497 5583 7531
rect 7941 7497 7975 7531
rect 4414 7429 4448 7463
rect 2717 7361 2751 7395
rect 6828 7361 6862 7395
rect 2973 7293 3007 7327
rect 4169 7293 4203 7327
rect 6561 7293 6595 7327
rect 3249 6817 3283 6851
rect 1777 6749 1811 6783
rect 2973 6749 3007 6783
rect 3433 6749 3467 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 4629 6749 4663 6783
rect 5457 6749 5491 6783
rect 3065 6681 3099 6715
rect 5724 6681 5758 6715
rect 1593 6613 1627 6647
rect 6837 6613 6871 6647
rect 4077 6409 4111 6443
rect 5825 6409 5859 6443
rect 6653 6409 6687 6443
rect 4261 6273 4295 6307
rect 4445 6273 4479 6307
rect 4537 6273 4571 6307
rect 5457 6273 5491 6307
rect 5641 6273 5675 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 5365 6205 5399 6239
rect 4445 5865 4479 5899
rect 5089 5865 5123 5899
rect 5273 5865 5307 5899
rect 6009 5865 6043 5899
rect 3433 5729 3467 5763
rect 4077 5729 4111 5763
rect 3157 5661 3191 5695
rect 3249 5661 3283 5695
rect 4261 5661 4295 5695
rect 5733 5661 5767 5695
rect 4905 5593 4939 5627
rect 5121 5593 5155 5627
rect 6009 5593 6043 5627
rect 3433 5525 3467 5559
rect 5825 5525 5859 5559
rect 2973 5321 3007 5355
rect 3985 5321 4019 5355
rect 7941 5321 7975 5355
rect 5917 5253 5951 5287
rect 3157 5185 3191 5219
rect 3341 5185 3375 5219
rect 4353 5185 4387 5219
rect 4997 5185 5031 5219
rect 5273 5185 5307 5219
rect 5733 5185 5767 5219
rect 6009 5185 6043 5219
rect 6817 5185 6851 5219
rect 6561 5117 6595 5151
rect 5733 5049 5767 5083
rect 3157 4981 3191 5015
rect 3801 4981 3835 5015
rect 3985 4981 4019 5015
rect 4813 4981 4847 5015
rect 5181 4981 5215 5015
rect 5825 4777 5859 4811
rect 6561 4777 6595 4811
rect 3433 4573 3467 4607
rect 4445 4573 4479 4607
rect 4712 4573 4746 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 1685 4505 1719 4539
rect 1869 4505 1903 4539
rect 3249 4437 3283 4471
rect 3240 4165 3274 4199
rect 2973 4097 3007 4131
rect 4353 3893 4387 3927
rect 7849 3077 7883 3111
rect 8033 3009 8067 3043
rect 1869 2397 1903 2431
rect 4261 2397 4295 2431
rect 7849 2397 7883 2431
rect 1685 2261 1719 2295
rect 4077 2261 4111 2295
rect 8033 2261 8067 2295
<< metal1 >>
rect 1104 9274 8648 9296
rect 1104 9222 1893 9274
rect 1945 9222 1957 9274
rect 2009 9222 2021 9274
rect 2073 9222 2085 9274
rect 2137 9222 2149 9274
rect 2201 9222 3779 9274
rect 3831 9222 3843 9274
rect 3895 9222 3907 9274
rect 3959 9222 3971 9274
rect 4023 9222 4035 9274
rect 4087 9222 5665 9274
rect 5717 9222 5729 9274
rect 5781 9222 5793 9274
rect 5845 9222 5857 9274
rect 5909 9222 5921 9274
rect 5973 9222 7551 9274
rect 7603 9222 7615 9274
rect 7667 9222 7679 9274
rect 7731 9222 7743 9274
rect 7795 9222 7807 9274
rect 7859 9222 8648 9274
rect 1104 9200 8648 9222
rect 1302 9120 1308 9172
rect 1360 9160 1366 9172
rect 1765 9163 1823 9169
rect 1765 9160 1777 9163
rect 1360 9132 1777 9160
rect 1360 9120 1366 9132
rect 1765 9129 1777 9132
rect 1811 9129 1823 9163
rect 1765 9123 1823 9129
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6236 9132 6745 9160
rect 6236 9120 6242 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 9398 9160 9404 9172
rect 8067 9132 9404 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1544 8928 1593 8956
rect 1544 8916 1550 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 5592 8928 6561 8956
rect 5592 8916 5598 8928
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8956 7895 8959
rect 8110 8956 8116 8968
rect 7883 8928 8116 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 1104 8730 8648 8752
rect 1104 8678 2553 8730
rect 2605 8678 2617 8730
rect 2669 8678 2681 8730
rect 2733 8678 2745 8730
rect 2797 8678 2809 8730
rect 2861 8678 4439 8730
rect 4491 8678 4503 8730
rect 4555 8678 4567 8730
rect 4619 8678 4631 8730
rect 4683 8678 4695 8730
rect 4747 8678 6325 8730
rect 6377 8678 6389 8730
rect 6441 8678 6453 8730
rect 6505 8678 6517 8730
rect 6569 8678 6581 8730
rect 6633 8678 8211 8730
rect 8263 8678 8275 8730
rect 8327 8678 8339 8730
rect 8391 8678 8403 8730
rect 8455 8678 8467 8730
rect 8519 8678 8648 8730
rect 1104 8656 8648 8678
rect 1762 8616 1768 8628
rect 1723 8588 1768 8616
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 1104 8186 8648 8208
rect 1104 8134 1893 8186
rect 1945 8134 1957 8186
rect 2009 8134 2021 8186
rect 2073 8134 2085 8186
rect 2137 8134 2149 8186
rect 2201 8134 3779 8186
rect 3831 8134 3843 8186
rect 3895 8134 3907 8186
rect 3959 8134 3971 8186
rect 4023 8134 4035 8186
rect 4087 8134 5665 8186
rect 5717 8134 5729 8186
rect 5781 8134 5793 8186
rect 5845 8134 5857 8186
rect 5909 8134 5921 8186
rect 5973 8134 7551 8186
rect 7603 8134 7615 8186
rect 7667 8134 7679 8186
rect 7731 8134 7743 8186
rect 7795 8134 7807 8186
rect 7859 8134 8648 8186
rect 1104 8112 8648 8134
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4396 7840 4445 7868
rect 4396 7828 4402 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4890 7868 4896 7880
rect 4851 7840 4896 7868
rect 4433 7831 4491 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5074 7868 5080 7880
rect 5035 7840 5080 7868
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 7926 7868 7932 7880
rect 7883 7840 7932 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 4246 7732 4252 7744
rect 4207 7704 4252 7732
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4982 7732 4988 7744
rect 4943 7704 4988 7732
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 8018 7732 8024 7744
rect 7979 7704 8024 7732
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 1104 7642 8648 7664
rect 1104 7590 2553 7642
rect 2605 7590 2617 7642
rect 2669 7590 2681 7642
rect 2733 7590 2745 7642
rect 2797 7590 2809 7642
rect 2861 7590 4439 7642
rect 4491 7590 4503 7642
rect 4555 7590 4567 7642
rect 4619 7590 4631 7642
rect 4683 7590 4695 7642
rect 4747 7590 6325 7642
rect 6377 7590 6389 7642
rect 6441 7590 6453 7642
rect 6505 7590 6517 7642
rect 6569 7590 6581 7642
rect 6633 7590 8211 7642
rect 8263 7590 8275 7642
rect 8327 7590 8339 7642
rect 8391 7590 8403 7642
rect 8455 7590 8467 7642
rect 8519 7590 8648 7642
rect 1104 7568 8648 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 5534 7528 5540 7540
rect 5495 7500 5540 7528
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 7926 7528 7932 7540
rect 7887 7500 7932 7528
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4402 7463 4460 7469
rect 4402 7460 4414 7463
rect 4304 7432 4414 7460
rect 4304 7420 4310 7432
rect 4402 7429 4414 7432
rect 4448 7429 4460 7463
rect 4402 7423 4460 7429
rect 2705 7395 2763 7401
rect 2705 7361 2717 7395
rect 2751 7392 2763 7395
rect 3234 7392 3240 7404
rect 2751 7364 3240 7392
rect 2751 7361 2763 7364
rect 2705 7355 2763 7361
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 6822 7401 6828 7404
rect 6816 7392 6828 7401
rect 6783 7364 6828 7392
rect 6816 7355 6828 7364
rect 6822 7352 6828 7355
rect 6880 7352 6886 7404
rect 2961 7327 3019 7333
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 3007 7296 4169 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 4157 7293 4169 7296
rect 4203 7293 4215 7327
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 4157 7287 4215 7293
rect 5460 7296 6561 7324
rect 4172 7188 4200 7287
rect 5460 7200 5488 7296
rect 6549 7293 6561 7296
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 5442 7188 5448 7200
rect 4172 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 1104 7098 8648 7120
rect 1104 7046 1893 7098
rect 1945 7046 1957 7098
rect 2009 7046 2021 7098
rect 2073 7046 2085 7098
rect 2137 7046 2149 7098
rect 2201 7046 3779 7098
rect 3831 7046 3843 7098
rect 3895 7046 3907 7098
rect 3959 7046 3971 7098
rect 4023 7046 4035 7098
rect 4087 7046 5665 7098
rect 5717 7046 5729 7098
rect 5781 7046 5793 7098
rect 5845 7046 5857 7098
rect 5909 7046 5921 7098
rect 5973 7046 7551 7098
rect 7603 7046 7615 7098
rect 7667 7046 7679 7098
rect 7731 7046 7743 7098
rect 7795 7046 7807 7098
rect 7859 7046 8648 7098
rect 1104 7024 8648 7046
rect 3234 6848 3240 6860
rect 3195 6820 3240 6848
rect 3234 6808 3240 6820
rect 3292 6808 3298 6860
rect 4062 6848 4068 6860
rect 3344 6820 4068 6848
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6780 3019 6783
rect 3344 6780 3372 6820
rect 4062 6808 4068 6820
rect 4120 6848 4126 6860
rect 4120 6820 4476 6848
rect 4120 6808 4126 6820
rect 3007 6752 3372 6780
rect 3421 6783 3479 6789
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3467 6752 3985 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 4154 6780 4160 6792
rect 4115 6752 4160 6780
rect 3973 6743 4031 6749
rect 1780 6712 1808 6743
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4448 6789 4476 6820
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 4617 6743 4675 6749
rect 3053 6715 3111 6721
rect 3053 6712 3065 6715
rect 1780 6684 3065 6712
rect 3053 6681 3065 6684
rect 3099 6712 3111 6715
rect 4632 6712 4660 6743
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 3099 6684 4660 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1544 6616 1593 6644
rect 1544 6604 1550 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 4632 6644 4660 6684
rect 5712 6715 5770 6721
rect 5712 6681 5724 6715
rect 5758 6712 5770 6715
rect 5810 6712 5816 6724
rect 5758 6684 5816 6712
rect 5758 6681 5770 6684
rect 5712 6675 5770 6681
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 4632 6616 6837 6644
rect 1581 6607 1639 6613
rect 6825 6613 6837 6616
rect 6871 6644 6883 6647
rect 7098 6644 7104 6656
rect 6871 6616 7104 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 1104 6554 8648 6576
rect 1104 6502 2553 6554
rect 2605 6502 2617 6554
rect 2669 6502 2681 6554
rect 2733 6502 2745 6554
rect 2797 6502 2809 6554
rect 2861 6502 4439 6554
rect 4491 6502 4503 6554
rect 4555 6502 4567 6554
rect 4619 6502 4631 6554
rect 4683 6502 4695 6554
rect 4747 6502 6325 6554
rect 6377 6502 6389 6554
rect 6441 6502 6453 6554
rect 6505 6502 6517 6554
rect 6569 6502 6581 6554
rect 6633 6502 8211 6554
rect 8263 6502 8275 6554
rect 8327 6502 8339 6554
rect 8391 6502 8403 6554
rect 8455 6502 8467 6554
rect 8519 6502 8648 6554
rect 1104 6480 8648 6502
rect 4062 6440 4068 6452
rect 4023 6412 4068 6440
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4890 6440 4896 6452
rect 4212 6412 4896 6440
rect 4212 6400 4218 6412
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5810 6440 5816 6452
rect 5771 6412 5816 6440
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6822 6440 6828 6452
rect 6687 6412 6828 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 5534 6372 5540 6384
rect 4264 6344 5540 6372
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 4264 6313 4292 6344
rect 5534 6332 5540 6344
rect 5592 6332 5598 6384
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 3476 6276 4261 6304
rect 3476 6264 3482 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4430 6304 4436 6316
rect 4391 6276 4436 6304
rect 4249 6267 4307 6273
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4580 6276 4625 6304
rect 4580 6264 4586 6276
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 5258 6304 5264 6316
rect 5132 6276 5264 6304
rect 5132 6264 5138 6276
rect 5258 6264 5264 6276
rect 5316 6304 5322 6316
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 5316 6276 5457 6304
rect 5316 6264 5322 6276
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 5994 6304 6000 6316
rect 5675 6276 6000 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6236 6276 6561 6304
rect 6236 6264 6242 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6205 5411 6239
rect 5353 6199 5411 6205
rect 5368 6168 5396 6199
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6748 6236 6776 6267
rect 6144 6208 6776 6236
rect 6144 6196 6150 6208
rect 7098 6168 7104 6180
rect 5368 6140 7104 6168
rect 7098 6128 7104 6140
rect 7156 6128 7162 6180
rect 1104 6010 8648 6032
rect 1104 5958 1893 6010
rect 1945 5958 1957 6010
rect 2009 5958 2021 6010
rect 2073 5958 2085 6010
rect 2137 5958 2149 6010
rect 2201 5958 3779 6010
rect 3831 5958 3843 6010
rect 3895 5958 3907 6010
rect 3959 5958 3971 6010
rect 4023 5958 4035 6010
rect 4087 5958 5665 6010
rect 5717 5958 5729 6010
rect 5781 5958 5793 6010
rect 5845 5958 5857 6010
rect 5909 5958 5921 6010
rect 5973 5958 7551 6010
rect 7603 5958 7615 6010
rect 7667 5958 7679 6010
rect 7731 5958 7743 6010
rect 7795 5958 7807 6010
rect 7859 5958 8648 6010
rect 1104 5936 8648 5958
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4396 5868 4445 5896
rect 4396 5856 4402 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 5077 5899 5135 5905
rect 5077 5865 5089 5899
rect 5123 5865 5135 5899
rect 5258 5896 5264 5908
rect 5219 5868 5264 5896
rect 5077 5859 5135 5865
rect 4522 5828 4528 5840
rect 3252 5800 4528 5828
rect 3252 5704 3280 5800
rect 4522 5788 4528 5800
rect 4580 5828 4586 5840
rect 5092 5828 5120 5859
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 5994 5896 6000 5908
rect 5955 5868 6000 5896
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 4580 5800 5120 5828
rect 4580 5788 4586 5800
rect 3418 5760 3424 5772
rect 3379 5732 3424 5760
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4154 5760 4160 5772
rect 4111 5732 4160 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 3142 5692 3148 5704
rect 3103 5664 3148 5692
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3234 5652 3240 5704
rect 3292 5692 3298 5704
rect 4249 5695 4307 5701
rect 3292 5664 3337 5692
rect 3292 5652 3298 5664
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4982 5692 4988 5704
rect 4295 5664 4988 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5258 5652 5264 5704
rect 5316 5692 5322 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5316 5664 5733 5692
rect 5316 5652 5322 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 3160 5624 3188 5652
rect 4430 5624 4436 5636
rect 3160 5596 4436 5624
rect 4430 5584 4436 5596
rect 4488 5624 4494 5636
rect 4893 5627 4951 5633
rect 4893 5624 4905 5627
rect 4488 5596 4905 5624
rect 4488 5584 4494 5596
rect 4893 5593 4905 5596
rect 4939 5593 4951 5627
rect 4893 5587 4951 5593
rect 5109 5627 5167 5633
rect 5109 5593 5121 5627
rect 5155 5624 5167 5627
rect 5534 5624 5540 5636
rect 5155 5596 5540 5624
rect 5155 5593 5167 5596
rect 5109 5587 5167 5593
rect 3421 5559 3479 5565
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 3970 5556 3976 5568
rect 3467 5528 3976 5556
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4908 5556 4936 5587
rect 5534 5584 5540 5596
rect 5592 5584 5598 5636
rect 5994 5624 6000 5636
rect 5955 5596 6000 5624
rect 5994 5584 6000 5596
rect 6052 5584 6058 5636
rect 5258 5556 5264 5568
rect 4908 5528 5264 5556
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 7098 5556 7104 5568
rect 5859 5528 7104 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 1104 5466 8648 5488
rect 1104 5414 2553 5466
rect 2605 5414 2617 5466
rect 2669 5414 2681 5466
rect 2733 5414 2745 5466
rect 2797 5414 2809 5466
rect 2861 5414 4439 5466
rect 4491 5414 4503 5466
rect 4555 5414 4567 5466
rect 4619 5414 4631 5466
rect 4683 5414 4695 5466
rect 4747 5414 6325 5466
rect 6377 5414 6389 5466
rect 6441 5414 6453 5466
rect 6505 5414 6517 5466
rect 6569 5414 6581 5466
rect 6633 5414 8211 5466
rect 8263 5414 8275 5466
rect 8327 5414 8339 5466
rect 8391 5414 8403 5466
rect 8455 5414 8467 5466
rect 8519 5414 8648 5466
rect 1104 5392 8648 5414
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 3973 5355 4031 5361
rect 3973 5352 3985 5355
rect 3007 5324 3985 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 3973 5321 3985 5324
rect 4019 5321 4031 5355
rect 4890 5352 4896 5364
rect 3973 5315 4031 5321
rect 4356 5324 4896 5352
rect 3142 5216 3148 5228
rect 3103 5188 3148 5216
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3418 5216 3424 5228
rect 3375 5188 3424 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 4356 5225 4384 5324
rect 4890 5312 4896 5324
rect 4948 5352 4954 5364
rect 5994 5352 6000 5364
rect 4948 5324 6000 5352
rect 4948 5312 4954 5324
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 7929 5355 7987 5361
rect 7929 5352 7941 5355
rect 6886 5324 7941 5352
rect 5905 5287 5963 5293
rect 5905 5284 5917 5287
rect 5276 5256 5917 5284
rect 5276 5228 5304 5256
rect 5905 5253 5917 5256
rect 5951 5284 5963 5287
rect 6886 5284 6914 5324
rect 7929 5321 7941 5324
rect 7975 5352 7987 5355
rect 8110 5352 8116 5364
rect 7975 5324 8116 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 5951 5256 6914 5284
rect 5951 5253 5963 5256
rect 5905 5247 5963 5253
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5031 5188 5212 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5184 5080 5212 5188
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 5721 5219 5779 5225
rect 5316 5188 5361 5216
rect 5316 5176 5322 5188
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5216 6055 5219
rect 6178 5216 6184 5228
rect 6043 5188 6184 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 5736 5148 5764 5179
rect 5902 5148 5908 5160
rect 5736 5120 5908 5148
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 5721 5083 5779 5089
rect 5721 5080 5733 5083
rect 3160 5052 4936 5080
rect 5184 5052 5733 5080
rect 3160 5024 3188 5052
rect 3142 5012 3148 5024
rect 3103 4984 3148 5012
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3476 4984 3801 5012
rect 3476 4972 3482 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 3970 5012 3976 5024
rect 3931 4984 3976 5012
rect 3789 4975 3847 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 4764 4984 4813 5012
rect 4764 4972 4770 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 4908 5012 4936 5052
rect 5721 5049 5733 5052
rect 5767 5049 5779 5083
rect 5721 5043 5779 5049
rect 5169 5015 5227 5021
rect 5169 5012 5181 5015
rect 4908 4984 5181 5012
rect 4801 4975 4859 4981
rect 5169 4981 5181 4984
rect 5215 5012 5227 5015
rect 5534 5012 5540 5024
rect 5215 4984 5540 5012
rect 5215 4981 5227 4984
rect 5169 4975 5227 4981
rect 5534 4972 5540 4984
rect 5592 5012 5598 5024
rect 6012 5012 6040 5179
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 6805 5219 6863 5225
rect 6805 5216 6817 5219
rect 6696 5188 6817 5216
rect 6696 5176 6702 5188
rect 6805 5185 6817 5188
rect 6851 5185 6863 5219
rect 6805 5179 6863 5185
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6549 5151 6607 5157
rect 6549 5148 6561 5151
rect 6512 5120 6561 5148
rect 6512 5108 6518 5120
rect 6549 5117 6561 5120
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 5592 4984 6040 5012
rect 5592 4972 5598 4984
rect 1104 4922 8648 4944
rect 1104 4870 1893 4922
rect 1945 4870 1957 4922
rect 2009 4870 2021 4922
rect 2073 4870 2085 4922
rect 2137 4870 2149 4922
rect 2201 4870 3779 4922
rect 3831 4870 3843 4922
rect 3895 4870 3907 4922
rect 3959 4870 3971 4922
rect 4023 4870 4035 4922
rect 4087 4870 5665 4922
rect 5717 4870 5729 4922
rect 5781 4870 5793 4922
rect 5845 4870 5857 4922
rect 5909 4870 5921 4922
rect 5973 4870 7551 4922
rect 7603 4870 7615 4922
rect 7667 4870 7679 4922
rect 7731 4870 7743 4922
rect 7795 4870 7807 4922
rect 7859 4870 8648 4922
rect 1104 4848 8648 4870
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5592 4780 5825 4808
rect 5592 4768 5598 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 6549 4811 6607 4817
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 6638 4808 6644 4820
rect 6595 4780 6644 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6052 4644 6592 4672
rect 6052 4632 6058 4644
rect 3418 4604 3424 4616
rect 3379 4576 3424 4604
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 4706 4613 4712 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4700 4604 4712 4613
rect 4667 4576 4712 4604
rect 4433 4567 4491 4573
rect 4700 4567 4712 4576
rect 1670 4536 1676 4548
rect 1631 4508 1676 4536
rect 1670 4496 1676 4508
rect 1728 4496 1734 4548
rect 1857 4539 1915 4545
rect 1857 4505 1869 4539
rect 1903 4536 1915 4539
rect 2958 4536 2964 4548
rect 1903 4508 2964 4536
rect 1903 4505 1915 4508
rect 1857 4499 1915 4505
rect 2958 4496 2964 4508
rect 3016 4536 3022 4548
rect 4448 4536 4476 4567
rect 4706 4564 4712 4567
rect 4764 4564 4770 4616
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 6564 4613 6592 4644
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 5316 4576 6377 4604
rect 5316 4564 5322 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4604 6607 4607
rect 6730 4604 6736 4616
rect 6595 4576 6736 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 5442 4536 5448 4548
rect 3016 4508 5448 4536
rect 3016 4496 3022 4508
rect 5442 4496 5448 4508
rect 5500 4536 5506 4548
rect 6454 4536 6460 4548
rect 5500 4508 6460 4536
rect 5500 4496 5506 4508
rect 6454 4496 6460 4508
rect 6512 4496 6518 4548
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 1104 4378 8648 4400
rect 1104 4326 2553 4378
rect 2605 4326 2617 4378
rect 2669 4326 2681 4378
rect 2733 4326 2745 4378
rect 2797 4326 2809 4378
rect 2861 4326 4439 4378
rect 4491 4326 4503 4378
rect 4555 4326 4567 4378
rect 4619 4326 4631 4378
rect 4683 4326 4695 4378
rect 4747 4326 6325 4378
rect 6377 4326 6389 4378
rect 6441 4326 6453 4378
rect 6505 4326 6517 4378
rect 6569 4326 6581 4378
rect 6633 4326 8211 4378
rect 8263 4326 8275 4378
rect 8327 4326 8339 4378
rect 8391 4326 8403 4378
rect 8455 4326 8467 4378
rect 8519 4326 8648 4378
rect 1104 4304 8648 4326
rect 3234 4205 3240 4208
rect 3228 4196 3240 4205
rect 3195 4168 3240 4196
rect 3228 4159 3240 4168
rect 3234 4156 3240 4159
rect 3292 4156 3298 4208
rect 2958 4128 2964 4140
rect 2919 4100 2964 4128
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 4304 3896 4353 3924
rect 4304 3884 4310 3896
rect 4341 3893 4353 3896
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 1104 3834 8648 3856
rect 1104 3782 1893 3834
rect 1945 3782 1957 3834
rect 2009 3782 2021 3834
rect 2073 3782 2085 3834
rect 2137 3782 2149 3834
rect 2201 3782 3779 3834
rect 3831 3782 3843 3834
rect 3895 3782 3907 3834
rect 3959 3782 3971 3834
rect 4023 3782 4035 3834
rect 4087 3782 5665 3834
rect 5717 3782 5729 3834
rect 5781 3782 5793 3834
rect 5845 3782 5857 3834
rect 5909 3782 5921 3834
rect 5973 3782 7551 3834
rect 7603 3782 7615 3834
rect 7667 3782 7679 3834
rect 7731 3782 7743 3834
rect 7795 3782 7807 3834
rect 7859 3782 8648 3834
rect 1104 3760 8648 3782
rect 1104 3290 8648 3312
rect 1104 3238 2553 3290
rect 2605 3238 2617 3290
rect 2669 3238 2681 3290
rect 2733 3238 2745 3290
rect 2797 3238 2809 3290
rect 2861 3238 4439 3290
rect 4491 3238 4503 3290
rect 4555 3238 4567 3290
rect 4619 3238 4631 3290
rect 4683 3238 4695 3290
rect 4747 3238 6325 3290
rect 6377 3238 6389 3290
rect 6441 3238 6453 3290
rect 6505 3238 6517 3290
rect 6569 3238 6581 3290
rect 6633 3238 8211 3290
rect 8263 3238 8275 3290
rect 8327 3238 8339 3290
rect 8391 3238 8403 3290
rect 8455 3238 8467 3290
rect 8519 3238 8648 3290
rect 1104 3216 8648 3238
rect 6730 3068 6736 3120
rect 6788 3108 6794 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 6788 3080 7849 3108
rect 6788 3068 6794 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 8018 3040 8024 3052
rect 7979 3012 8024 3040
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 1104 2746 8648 2768
rect 1104 2694 1893 2746
rect 1945 2694 1957 2746
rect 2009 2694 2021 2746
rect 2073 2694 2085 2746
rect 2137 2694 2149 2746
rect 2201 2694 3779 2746
rect 3831 2694 3843 2746
rect 3895 2694 3907 2746
rect 3959 2694 3971 2746
rect 4023 2694 4035 2746
rect 4087 2694 5665 2746
rect 5717 2694 5729 2746
rect 5781 2694 5793 2746
rect 5845 2694 5857 2746
rect 5909 2694 5921 2746
rect 5973 2694 7551 2746
rect 7603 2694 7615 2746
rect 7667 2694 7679 2746
rect 7731 2694 7743 2746
rect 7795 2694 7807 2746
rect 7859 2694 8648 2746
rect 1104 2672 8648 2694
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 3142 2428 3148 2440
rect 1903 2400 3148 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 4246 2428 4252 2440
rect 4207 2400 4252 2428
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7156 2400 7849 2428
rect 7156 2388 7162 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 72 2264 1685 2292
rect 72 2252 78 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 8021 2295 8079 2301
rect 8021 2261 8033 2295
rect 8067 2292 8079 2295
rect 8110 2292 8116 2304
rect 8067 2264 8116 2292
rect 8067 2261 8079 2264
rect 8021 2255 8079 2261
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 1104 2202 8648 2224
rect 1104 2150 2553 2202
rect 2605 2150 2617 2202
rect 2669 2150 2681 2202
rect 2733 2150 2745 2202
rect 2797 2150 2809 2202
rect 2861 2150 4439 2202
rect 4491 2150 4503 2202
rect 4555 2150 4567 2202
rect 4619 2150 4631 2202
rect 4683 2150 4695 2202
rect 4747 2150 6325 2202
rect 6377 2150 6389 2202
rect 6441 2150 6453 2202
rect 6505 2150 6517 2202
rect 6569 2150 6581 2202
rect 6633 2150 8211 2202
rect 8263 2150 8275 2202
rect 8327 2150 8339 2202
rect 8391 2150 8403 2202
rect 8455 2150 8467 2202
rect 8519 2150 8648 2202
rect 1104 2128 8648 2150
<< via1 >>
rect 1893 9222 1945 9274
rect 1957 9222 2009 9274
rect 2021 9222 2073 9274
rect 2085 9222 2137 9274
rect 2149 9222 2201 9274
rect 3779 9222 3831 9274
rect 3843 9222 3895 9274
rect 3907 9222 3959 9274
rect 3971 9222 4023 9274
rect 4035 9222 4087 9274
rect 5665 9222 5717 9274
rect 5729 9222 5781 9274
rect 5793 9222 5845 9274
rect 5857 9222 5909 9274
rect 5921 9222 5973 9274
rect 7551 9222 7603 9274
rect 7615 9222 7667 9274
rect 7679 9222 7731 9274
rect 7743 9222 7795 9274
rect 7807 9222 7859 9274
rect 1308 9120 1360 9172
rect 6184 9120 6236 9172
rect 9404 9120 9456 9172
rect 1492 8916 1544 8968
rect 5540 8916 5592 8968
rect 8116 8916 8168 8968
rect 2553 8678 2605 8730
rect 2617 8678 2669 8730
rect 2681 8678 2733 8730
rect 2745 8678 2797 8730
rect 2809 8678 2861 8730
rect 4439 8678 4491 8730
rect 4503 8678 4555 8730
rect 4567 8678 4619 8730
rect 4631 8678 4683 8730
rect 4695 8678 4747 8730
rect 6325 8678 6377 8730
rect 6389 8678 6441 8730
rect 6453 8678 6505 8730
rect 6517 8678 6569 8730
rect 6581 8678 6633 8730
rect 8211 8678 8263 8730
rect 8275 8678 8327 8730
rect 8339 8678 8391 8730
rect 8403 8678 8455 8730
rect 8467 8678 8519 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 1893 8134 1945 8186
rect 1957 8134 2009 8186
rect 2021 8134 2073 8186
rect 2085 8134 2137 8186
rect 2149 8134 2201 8186
rect 3779 8134 3831 8186
rect 3843 8134 3895 8186
rect 3907 8134 3959 8186
rect 3971 8134 4023 8186
rect 4035 8134 4087 8186
rect 5665 8134 5717 8186
rect 5729 8134 5781 8186
rect 5793 8134 5845 8186
rect 5857 8134 5909 8186
rect 5921 8134 5973 8186
rect 7551 8134 7603 8186
rect 7615 8134 7667 8186
rect 7679 8134 7731 8186
rect 7743 8134 7795 8186
rect 7807 8134 7859 8186
rect 4344 7828 4396 7880
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 7932 7828 7984 7880
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 4988 7735 5040 7744
rect 4988 7701 4997 7735
rect 4997 7701 5031 7735
rect 5031 7701 5040 7735
rect 4988 7692 5040 7701
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 2553 7590 2605 7642
rect 2617 7590 2669 7642
rect 2681 7590 2733 7642
rect 2745 7590 2797 7642
rect 2809 7590 2861 7642
rect 4439 7590 4491 7642
rect 4503 7590 4555 7642
rect 4567 7590 4619 7642
rect 4631 7590 4683 7642
rect 4695 7590 4747 7642
rect 6325 7590 6377 7642
rect 6389 7590 6441 7642
rect 6453 7590 6505 7642
rect 6517 7590 6569 7642
rect 6581 7590 6633 7642
rect 8211 7590 8263 7642
rect 8275 7590 8327 7642
rect 8339 7590 8391 7642
rect 8403 7590 8455 7642
rect 8467 7590 8519 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 4252 7420 4304 7472
rect 3240 7352 3292 7404
rect 6828 7395 6880 7404
rect 6828 7361 6862 7395
rect 6862 7361 6880 7395
rect 6828 7352 6880 7361
rect 5448 7148 5500 7200
rect 1893 7046 1945 7098
rect 1957 7046 2009 7098
rect 2021 7046 2073 7098
rect 2085 7046 2137 7098
rect 2149 7046 2201 7098
rect 3779 7046 3831 7098
rect 3843 7046 3895 7098
rect 3907 7046 3959 7098
rect 3971 7046 4023 7098
rect 4035 7046 4087 7098
rect 5665 7046 5717 7098
rect 5729 7046 5781 7098
rect 5793 7046 5845 7098
rect 5857 7046 5909 7098
rect 5921 7046 5973 7098
rect 7551 7046 7603 7098
rect 7615 7046 7667 7098
rect 7679 7046 7731 7098
rect 7743 7046 7795 7098
rect 7807 7046 7859 7098
rect 3240 6851 3292 6860
rect 3240 6817 3249 6851
rect 3249 6817 3283 6851
rect 3283 6817 3292 6851
rect 3240 6808 3292 6817
rect 4068 6808 4120 6860
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 1492 6604 1544 6656
rect 5816 6672 5868 6724
rect 7104 6604 7156 6656
rect 2553 6502 2605 6554
rect 2617 6502 2669 6554
rect 2681 6502 2733 6554
rect 2745 6502 2797 6554
rect 2809 6502 2861 6554
rect 4439 6502 4491 6554
rect 4503 6502 4555 6554
rect 4567 6502 4619 6554
rect 4631 6502 4683 6554
rect 4695 6502 4747 6554
rect 6325 6502 6377 6554
rect 6389 6502 6441 6554
rect 6453 6502 6505 6554
rect 6517 6502 6569 6554
rect 6581 6502 6633 6554
rect 8211 6502 8263 6554
rect 8275 6502 8327 6554
rect 8339 6502 8391 6554
rect 8403 6502 8455 6554
rect 8467 6502 8519 6554
rect 4068 6443 4120 6452
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 4160 6400 4212 6452
rect 4896 6400 4948 6452
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 6828 6400 6880 6452
rect 3424 6264 3476 6316
rect 5540 6332 5592 6384
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 5080 6264 5132 6316
rect 5264 6264 5316 6316
rect 6000 6264 6052 6316
rect 6184 6264 6236 6316
rect 6092 6196 6144 6248
rect 7104 6128 7156 6180
rect 1893 5958 1945 6010
rect 1957 5958 2009 6010
rect 2021 5958 2073 6010
rect 2085 5958 2137 6010
rect 2149 5958 2201 6010
rect 3779 5958 3831 6010
rect 3843 5958 3895 6010
rect 3907 5958 3959 6010
rect 3971 5958 4023 6010
rect 4035 5958 4087 6010
rect 5665 5958 5717 6010
rect 5729 5958 5781 6010
rect 5793 5958 5845 6010
rect 5857 5958 5909 6010
rect 5921 5958 5973 6010
rect 7551 5958 7603 6010
rect 7615 5958 7667 6010
rect 7679 5958 7731 6010
rect 7743 5958 7795 6010
rect 7807 5958 7859 6010
rect 4344 5856 4396 5908
rect 5264 5899 5316 5908
rect 4528 5788 4580 5840
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 5264 5856 5316 5865
rect 6000 5899 6052 5908
rect 6000 5865 6009 5899
rect 6009 5865 6043 5899
rect 6043 5865 6052 5899
rect 6000 5856 6052 5865
rect 3424 5763 3476 5772
rect 3424 5729 3433 5763
rect 3433 5729 3467 5763
rect 3467 5729 3476 5763
rect 3424 5720 3476 5729
rect 4160 5720 4212 5772
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 4988 5652 5040 5704
rect 5264 5652 5316 5704
rect 4436 5584 4488 5636
rect 3976 5516 4028 5568
rect 5540 5584 5592 5636
rect 6000 5627 6052 5636
rect 6000 5593 6009 5627
rect 6009 5593 6043 5627
rect 6043 5593 6052 5627
rect 6000 5584 6052 5593
rect 5264 5516 5316 5568
rect 7104 5516 7156 5568
rect 2553 5414 2605 5466
rect 2617 5414 2669 5466
rect 2681 5414 2733 5466
rect 2745 5414 2797 5466
rect 2809 5414 2861 5466
rect 4439 5414 4491 5466
rect 4503 5414 4555 5466
rect 4567 5414 4619 5466
rect 4631 5414 4683 5466
rect 4695 5414 4747 5466
rect 6325 5414 6377 5466
rect 6389 5414 6441 5466
rect 6453 5414 6505 5466
rect 6517 5414 6569 5466
rect 6581 5414 6633 5466
rect 8211 5414 8263 5466
rect 8275 5414 8327 5466
rect 8339 5414 8391 5466
rect 8403 5414 8455 5466
rect 8467 5414 8519 5466
rect 3148 5219 3200 5228
rect 3148 5185 3157 5219
rect 3157 5185 3191 5219
rect 3191 5185 3200 5219
rect 3148 5176 3200 5185
rect 3424 5176 3476 5228
rect 4896 5312 4948 5364
rect 6000 5312 6052 5364
rect 8116 5312 8168 5364
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 5908 5108 5960 5160
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 3148 4972 3200 4981
rect 3424 4972 3476 5024
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 4712 4972 4764 5024
rect 5540 4972 5592 5024
rect 6184 5176 6236 5228
rect 6644 5176 6696 5228
rect 6460 5108 6512 5160
rect 1893 4870 1945 4922
rect 1957 4870 2009 4922
rect 2021 4870 2073 4922
rect 2085 4870 2137 4922
rect 2149 4870 2201 4922
rect 3779 4870 3831 4922
rect 3843 4870 3895 4922
rect 3907 4870 3959 4922
rect 3971 4870 4023 4922
rect 4035 4870 4087 4922
rect 5665 4870 5717 4922
rect 5729 4870 5781 4922
rect 5793 4870 5845 4922
rect 5857 4870 5909 4922
rect 5921 4870 5973 4922
rect 7551 4870 7603 4922
rect 7615 4870 7667 4922
rect 7679 4870 7731 4922
rect 7743 4870 7795 4922
rect 7807 4870 7859 4922
rect 5540 4768 5592 4820
rect 6644 4768 6696 4820
rect 6000 4632 6052 4684
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 4712 4607 4764 4616
rect 4712 4573 4746 4607
rect 4746 4573 4764 4607
rect 1676 4539 1728 4548
rect 1676 4505 1685 4539
rect 1685 4505 1719 4539
rect 1719 4505 1728 4539
rect 1676 4496 1728 4505
rect 2964 4496 3016 4548
rect 4712 4564 4764 4573
rect 5264 4564 5316 4616
rect 6736 4564 6788 4616
rect 5448 4496 5500 4548
rect 6460 4496 6512 4548
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 2553 4326 2605 4378
rect 2617 4326 2669 4378
rect 2681 4326 2733 4378
rect 2745 4326 2797 4378
rect 2809 4326 2861 4378
rect 4439 4326 4491 4378
rect 4503 4326 4555 4378
rect 4567 4326 4619 4378
rect 4631 4326 4683 4378
rect 4695 4326 4747 4378
rect 6325 4326 6377 4378
rect 6389 4326 6441 4378
rect 6453 4326 6505 4378
rect 6517 4326 6569 4378
rect 6581 4326 6633 4378
rect 8211 4326 8263 4378
rect 8275 4326 8327 4378
rect 8339 4326 8391 4378
rect 8403 4326 8455 4378
rect 8467 4326 8519 4378
rect 3240 4199 3292 4208
rect 3240 4165 3274 4199
rect 3274 4165 3292 4199
rect 3240 4156 3292 4165
rect 2964 4131 3016 4140
rect 2964 4097 2973 4131
rect 2973 4097 3007 4131
rect 3007 4097 3016 4131
rect 2964 4088 3016 4097
rect 4252 3884 4304 3936
rect 1893 3782 1945 3834
rect 1957 3782 2009 3834
rect 2021 3782 2073 3834
rect 2085 3782 2137 3834
rect 2149 3782 2201 3834
rect 3779 3782 3831 3834
rect 3843 3782 3895 3834
rect 3907 3782 3959 3834
rect 3971 3782 4023 3834
rect 4035 3782 4087 3834
rect 5665 3782 5717 3834
rect 5729 3782 5781 3834
rect 5793 3782 5845 3834
rect 5857 3782 5909 3834
rect 5921 3782 5973 3834
rect 7551 3782 7603 3834
rect 7615 3782 7667 3834
rect 7679 3782 7731 3834
rect 7743 3782 7795 3834
rect 7807 3782 7859 3834
rect 2553 3238 2605 3290
rect 2617 3238 2669 3290
rect 2681 3238 2733 3290
rect 2745 3238 2797 3290
rect 2809 3238 2861 3290
rect 4439 3238 4491 3290
rect 4503 3238 4555 3290
rect 4567 3238 4619 3290
rect 4631 3238 4683 3290
rect 4695 3238 4747 3290
rect 6325 3238 6377 3290
rect 6389 3238 6441 3290
rect 6453 3238 6505 3290
rect 6517 3238 6569 3290
rect 6581 3238 6633 3290
rect 8211 3238 8263 3290
rect 8275 3238 8327 3290
rect 8339 3238 8391 3290
rect 8403 3238 8455 3290
rect 8467 3238 8519 3290
rect 6736 3068 6788 3120
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 1893 2694 1945 2746
rect 1957 2694 2009 2746
rect 2021 2694 2073 2746
rect 2085 2694 2137 2746
rect 2149 2694 2201 2746
rect 3779 2694 3831 2746
rect 3843 2694 3895 2746
rect 3907 2694 3959 2746
rect 3971 2694 4023 2746
rect 4035 2694 4087 2746
rect 5665 2694 5717 2746
rect 5729 2694 5781 2746
rect 5793 2694 5845 2746
rect 5857 2694 5909 2746
rect 5921 2694 5973 2746
rect 7551 2694 7603 2746
rect 7615 2694 7667 2746
rect 7679 2694 7731 2746
rect 7743 2694 7795 2746
rect 7807 2694 7859 2746
rect 3148 2388 3200 2440
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 7104 2388 7156 2440
rect 20 2252 72 2304
rect 3884 2252 3936 2304
rect 8116 2252 8168 2304
rect 2553 2150 2605 2202
rect 2617 2150 2669 2202
rect 2681 2150 2733 2202
rect 2745 2150 2797 2202
rect 2809 2150 2861 2202
rect 4439 2150 4491 2202
rect 4503 2150 4555 2202
rect 4567 2150 4619 2202
rect 4631 2150 4683 2202
rect 4695 2150 4747 2202
rect 6325 2150 6377 2202
rect 6389 2150 6441 2202
rect 6453 2150 6505 2202
rect 6517 2150 6569 2202
rect 6581 2150 6633 2202
rect 8211 2150 8263 2202
rect 8275 2150 8327 2202
rect 8339 2150 8391 2202
rect 8403 2150 8455 2202
rect 8467 2150 8519 2202
<< metal2 >>
rect 1306 11122 1362 11922
rect 5814 11234 5870 11922
rect 9678 11234 9734 11922
rect 5814 11206 6224 11234
rect 5814 11122 5870 11206
rect 1320 9178 1348 11122
rect 1893 9276 2201 9285
rect 1893 9274 1899 9276
rect 1955 9274 1979 9276
rect 2035 9274 2059 9276
rect 2115 9274 2139 9276
rect 2195 9274 2201 9276
rect 1955 9222 1957 9274
rect 2137 9222 2139 9274
rect 1893 9220 1899 9222
rect 1955 9220 1979 9222
rect 2035 9220 2059 9222
rect 2115 9220 2139 9222
rect 2195 9220 2201 9222
rect 1893 9211 2201 9220
rect 3779 9276 4087 9285
rect 3779 9274 3785 9276
rect 3841 9274 3865 9276
rect 3921 9274 3945 9276
rect 4001 9274 4025 9276
rect 4081 9274 4087 9276
rect 3841 9222 3843 9274
rect 4023 9222 4025 9274
rect 3779 9220 3785 9222
rect 3841 9220 3865 9222
rect 3921 9220 3945 9222
rect 4001 9220 4025 9222
rect 4081 9220 4087 9222
rect 3779 9211 4087 9220
rect 5665 9276 5973 9285
rect 5665 9274 5671 9276
rect 5727 9274 5751 9276
rect 5807 9274 5831 9276
rect 5887 9274 5911 9276
rect 5967 9274 5973 9276
rect 5727 9222 5729 9274
rect 5909 9222 5911 9274
rect 5665 9220 5671 9222
rect 5727 9220 5751 9222
rect 5807 9220 5831 9222
rect 5887 9220 5911 9222
rect 5967 9220 5973 9222
rect 5665 9211 5973 9220
rect 6196 9178 6224 11206
rect 9416 11206 9734 11234
rect 7551 9276 7859 9285
rect 7551 9274 7557 9276
rect 7613 9274 7637 9276
rect 7693 9274 7717 9276
rect 7773 9274 7797 9276
rect 7853 9274 7859 9276
rect 7613 9222 7615 9274
rect 7795 9222 7797 9274
rect 7551 9220 7557 9222
rect 7613 9220 7637 9222
rect 7693 9220 7717 9222
rect 7773 9220 7797 9222
rect 7853 9220 7859 9222
rect 7551 9211 7859 9220
rect 9416 9178 9444 11206
rect 9678 11122 9734 11206
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 1492 8968 1544 8974
rect 5540 8968 5592 8974
rect 1492 8910 1544 8916
rect 1766 8936 1822 8945
rect 1504 6662 1532 8910
rect 5540 8910 5592 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 1766 8871 1822 8880
rect 1780 8634 1808 8871
rect 2553 8732 2861 8741
rect 2553 8730 2559 8732
rect 2615 8730 2639 8732
rect 2695 8730 2719 8732
rect 2775 8730 2799 8732
rect 2855 8730 2861 8732
rect 2615 8678 2617 8730
rect 2797 8678 2799 8730
rect 2553 8676 2559 8678
rect 2615 8676 2639 8678
rect 2695 8676 2719 8678
rect 2775 8676 2799 8678
rect 2855 8676 2861 8678
rect 2553 8667 2861 8676
rect 4439 8732 4747 8741
rect 4439 8730 4445 8732
rect 4501 8730 4525 8732
rect 4581 8730 4605 8732
rect 4661 8730 4685 8732
rect 4741 8730 4747 8732
rect 4501 8678 4503 8730
rect 4683 8678 4685 8730
rect 4439 8676 4445 8678
rect 4501 8676 4525 8678
rect 4581 8676 4605 8678
rect 4661 8676 4685 8678
rect 4741 8676 4747 8678
rect 4439 8667 4747 8676
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 7546 1624 8434
rect 1893 8188 2201 8197
rect 1893 8186 1899 8188
rect 1955 8186 1979 8188
rect 2035 8186 2059 8188
rect 2115 8186 2139 8188
rect 2195 8186 2201 8188
rect 1955 8134 1957 8186
rect 2137 8134 2139 8186
rect 1893 8132 1899 8134
rect 1955 8132 1979 8134
rect 2035 8132 2059 8134
rect 2115 8132 2139 8134
rect 2195 8132 2201 8134
rect 1893 8123 2201 8132
rect 3779 8188 4087 8197
rect 3779 8186 3785 8188
rect 3841 8186 3865 8188
rect 3921 8186 3945 8188
rect 4001 8186 4025 8188
rect 4081 8186 4087 8188
rect 3841 8134 3843 8186
rect 4023 8134 4025 8186
rect 3779 8132 3785 8134
rect 3841 8132 3865 8134
rect 3921 8132 3945 8134
rect 4001 8132 4025 8134
rect 4081 8132 4087 8134
rect 3779 8123 4087 8132
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 2553 7644 2861 7653
rect 2553 7642 2559 7644
rect 2615 7642 2639 7644
rect 2695 7642 2719 7644
rect 2775 7642 2799 7644
rect 2855 7642 2861 7644
rect 2615 7590 2617 7642
rect 2797 7590 2799 7642
rect 2553 7588 2559 7590
rect 2615 7588 2639 7590
rect 2695 7588 2719 7590
rect 2775 7588 2799 7590
rect 2855 7588 2861 7590
rect 2553 7579 2861 7588
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 4264 7478 4292 7686
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 1893 7100 2201 7109
rect 1893 7098 1899 7100
rect 1955 7098 1979 7100
rect 2035 7098 2059 7100
rect 2115 7098 2139 7100
rect 2195 7098 2201 7100
rect 1955 7046 1957 7098
rect 2137 7046 2139 7098
rect 1893 7044 1899 7046
rect 1955 7044 1979 7046
rect 2035 7044 2059 7046
rect 2115 7044 2139 7046
rect 2195 7044 2201 7046
rect 1893 7035 2201 7044
rect 3252 6866 3280 7346
rect 3779 7100 4087 7109
rect 3779 7098 3785 7100
rect 3841 7098 3865 7100
rect 3921 7098 3945 7100
rect 4001 7098 4025 7100
rect 4081 7098 4087 7100
rect 3841 7046 3843 7098
rect 4023 7046 4025 7098
rect 3779 7044 3785 7046
rect 3841 7044 3865 7046
rect 3921 7044 3945 7046
rect 4001 7044 4025 7046
rect 4081 7044 4087 7046
rect 3779 7035 4087 7044
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 2553 6556 2861 6565
rect 2553 6554 2559 6556
rect 2615 6554 2639 6556
rect 2695 6554 2719 6556
rect 2775 6554 2799 6556
rect 2855 6554 2861 6556
rect 2615 6502 2617 6554
rect 2797 6502 2799 6554
rect 2553 6500 2559 6502
rect 2615 6500 2639 6502
rect 2695 6500 2719 6502
rect 2775 6500 2799 6502
rect 2855 6500 2861 6502
rect 2553 6491 2861 6500
rect 4080 6458 4108 6802
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4172 6458 4200 6734
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 1893 6012 2201 6021
rect 1893 6010 1899 6012
rect 1955 6010 1979 6012
rect 2035 6010 2059 6012
rect 2115 6010 2139 6012
rect 2195 6010 2201 6012
rect 1955 5958 1957 6010
rect 2137 5958 2139 6010
rect 1893 5956 1899 5958
rect 1955 5956 1979 5958
rect 2035 5956 2059 5958
rect 2115 5956 2139 5958
rect 2195 5956 2201 5958
rect 1893 5947 2201 5956
rect 3436 5778 3464 6258
rect 4080 6202 4108 6394
rect 4080 6174 4200 6202
rect 3779 6012 4087 6021
rect 3779 6010 3785 6012
rect 3841 6010 3865 6012
rect 3921 6010 3945 6012
rect 4001 6010 4025 6012
rect 4081 6010 4087 6012
rect 3841 5958 3843 6010
rect 4023 5958 4025 6010
rect 3779 5956 3785 5958
rect 3841 5956 3865 5958
rect 3921 5956 3945 5958
rect 4001 5956 4025 5958
rect 4081 5956 4087 5958
rect 3779 5947 4087 5956
rect 4172 5778 4200 6174
rect 4356 5914 4384 7822
rect 4439 7644 4747 7653
rect 4439 7642 4445 7644
rect 4501 7642 4525 7644
rect 4581 7642 4605 7644
rect 4661 7642 4685 7644
rect 4741 7642 4747 7644
rect 4501 7590 4503 7642
rect 4683 7590 4685 7642
rect 4439 7588 4445 7590
rect 4501 7588 4525 7590
rect 4581 7588 4605 7590
rect 4661 7588 4685 7590
rect 4741 7588 4747 7590
rect 4439 7579 4747 7588
rect 4439 6556 4747 6565
rect 4439 6554 4445 6556
rect 4501 6554 4525 6556
rect 4581 6554 4605 6556
rect 4661 6554 4685 6556
rect 4741 6554 4747 6556
rect 4501 6502 4503 6554
rect 4683 6502 4685 6554
rect 4439 6500 4445 6502
rect 4501 6500 4525 6502
rect 4581 6500 4605 6502
rect 4661 6500 4685 6502
rect 4741 6500 4747 6502
rect 4439 6491 4747 6500
rect 4908 6458 4936 7822
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 2553 5468 2861 5477
rect 2553 5466 2559 5468
rect 2615 5466 2639 5468
rect 2695 5466 2719 5468
rect 2775 5466 2799 5468
rect 2855 5466 2861 5468
rect 2615 5414 2617 5466
rect 2797 5414 2799 5466
rect 2553 5412 2559 5414
rect 2615 5412 2639 5414
rect 2695 5412 2719 5414
rect 2775 5412 2799 5414
rect 2855 5412 2861 5414
rect 2553 5403 2861 5412
rect 3160 5234 3188 5646
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3252 5114 3280 5646
rect 3436 5234 3464 5714
rect 4448 5642 4476 6258
rect 4540 5846 4568 6258
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3160 5086 3280 5114
rect 3160 5030 3188 5086
rect 3988 5030 4016 5510
rect 4439 5468 4747 5477
rect 4439 5466 4445 5468
rect 4501 5466 4525 5468
rect 4581 5466 4605 5468
rect 4661 5466 4685 5468
rect 4741 5466 4747 5468
rect 4501 5414 4503 5466
rect 4683 5414 4685 5466
rect 4439 5412 4445 5414
rect 4501 5412 4525 5414
rect 4581 5412 4605 5414
rect 4661 5412 4685 5414
rect 4741 5412 4747 5414
rect 4439 5403 4747 5412
rect 4908 5370 4936 6394
rect 5000 5710 5028 7686
rect 5092 6322 5120 7822
rect 5552 7546 5580 8910
rect 6325 8732 6633 8741
rect 6325 8730 6331 8732
rect 6387 8730 6411 8732
rect 6467 8730 6491 8732
rect 6547 8730 6571 8732
rect 6627 8730 6633 8732
rect 6387 8678 6389 8730
rect 6569 8678 6571 8730
rect 6325 8676 6331 8678
rect 6387 8676 6411 8678
rect 6467 8676 6491 8678
rect 6547 8676 6571 8678
rect 6627 8676 6633 8678
rect 6325 8667 6633 8676
rect 5665 8188 5973 8197
rect 5665 8186 5671 8188
rect 5727 8186 5751 8188
rect 5807 8186 5831 8188
rect 5887 8186 5911 8188
rect 5967 8186 5973 8188
rect 5727 8134 5729 8186
rect 5909 8134 5911 8186
rect 5665 8132 5671 8134
rect 5727 8132 5751 8134
rect 5807 8132 5831 8134
rect 5887 8132 5911 8134
rect 5967 8132 5973 8134
rect 5665 8123 5973 8132
rect 7551 8188 7859 8197
rect 7551 8186 7557 8188
rect 7613 8186 7637 8188
rect 7693 8186 7717 8188
rect 7773 8186 7797 8188
rect 7853 8186 7859 8188
rect 7613 8134 7615 8186
rect 7795 8134 7797 8186
rect 7551 8132 7557 8134
rect 7613 8132 7637 8134
rect 7693 8132 7717 8134
rect 7773 8132 7797 8134
rect 7853 8132 7859 8134
rect 7551 8123 7859 8132
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 6325 7644 6633 7653
rect 6325 7642 6331 7644
rect 6387 7642 6411 7644
rect 6467 7642 6491 7644
rect 6547 7642 6571 7644
rect 6627 7642 6633 7644
rect 6387 7590 6389 7642
rect 6569 7590 6571 7642
rect 6325 7588 6331 7590
rect 6387 7588 6411 7590
rect 6467 7588 6491 7590
rect 6547 7588 6571 7590
rect 6627 7588 6633 7590
rect 6325 7579 6633 7588
rect 7944 7546 7972 7822
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6798 5488 7142
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 5914 5304 6258
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5276 5710 5304 5850
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 5276 5234 5304 5510
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 1893 4924 2201 4933
rect 1893 4922 1899 4924
rect 1955 4922 1979 4924
rect 2035 4922 2059 4924
rect 2115 4922 2139 4924
rect 2195 4922 2201 4924
rect 1955 4870 1957 4922
rect 2137 4870 2139 4922
rect 1893 4868 1899 4870
rect 1955 4868 1979 4870
rect 2035 4868 2059 4870
rect 2115 4868 2139 4870
rect 2195 4868 2201 4870
rect 1893 4859 2201 4868
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 1688 4185 1716 4490
rect 2553 4380 2861 4389
rect 2553 4378 2559 4380
rect 2615 4378 2639 4380
rect 2695 4378 2719 4380
rect 2775 4378 2799 4380
rect 2855 4378 2861 4380
rect 2615 4326 2617 4378
rect 2797 4326 2799 4378
rect 2553 4324 2559 4326
rect 2615 4324 2639 4326
rect 2695 4324 2719 4326
rect 2775 4324 2799 4326
rect 2855 4324 2861 4326
rect 2553 4315 2861 4324
rect 1674 4176 1730 4185
rect 2976 4146 3004 4490
rect 1674 4111 1730 4120
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 1893 3836 2201 3845
rect 1893 3834 1899 3836
rect 1955 3834 1979 3836
rect 2035 3834 2059 3836
rect 2115 3834 2139 3836
rect 2195 3834 2201 3836
rect 1955 3782 1957 3834
rect 2137 3782 2139 3834
rect 1893 3780 1899 3782
rect 1955 3780 1979 3782
rect 2035 3780 2059 3782
rect 2115 3780 2139 3782
rect 2195 3780 2201 3782
rect 1893 3771 2201 3780
rect 2553 3292 2861 3301
rect 2553 3290 2559 3292
rect 2615 3290 2639 3292
rect 2695 3290 2719 3292
rect 2775 3290 2799 3292
rect 2855 3290 2861 3292
rect 2615 3238 2617 3290
rect 2797 3238 2799 3290
rect 2553 3236 2559 3238
rect 2615 3236 2639 3238
rect 2695 3236 2719 3238
rect 2775 3236 2799 3238
rect 2855 3236 2861 3238
rect 2553 3227 2861 3236
rect 1893 2748 2201 2757
rect 1893 2746 1899 2748
rect 1955 2746 1979 2748
rect 2035 2746 2059 2748
rect 2115 2746 2139 2748
rect 2195 2746 2201 2748
rect 1955 2694 1957 2746
rect 2137 2694 2139 2746
rect 1893 2692 1899 2694
rect 1955 2692 1979 2694
rect 2035 2692 2059 2694
rect 2115 2692 2139 2694
rect 2195 2692 2201 2694
rect 1893 2683 2201 2692
rect 3160 2446 3188 4966
rect 3436 4622 3464 4966
rect 3779 4924 4087 4933
rect 3779 4922 3785 4924
rect 3841 4922 3865 4924
rect 3921 4922 3945 4924
rect 4001 4922 4025 4924
rect 4081 4922 4087 4924
rect 3841 4870 3843 4922
rect 4023 4870 4025 4922
rect 3779 4868 3785 4870
rect 3841 4868 3865 4870
rect 3921 4868 3945 4870
rect 4001 4868 4025 4870
rect 4081 4868 4087 4870
rect 3779 4859 4087 4868
rect 4724 4622 4752 4966
rect 5276 4622 5304 5170
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5460 4554 5488 6734
rect 5552 6390 5580 7482
rect 8036 7449 8064 7686
rect 8022 7440 8078 7449
rect 6828 7404 6880 7410
rect 8022 7375 8078 7384
rect 6828 7346 6880 7352
rect 5665 7100 5973 7109
rect 5665 7098 5671 7100
rect 5727 7098 5751 7100
rect 5807 7098 5831 7100
rect 5887 7098 5911 7100
rect 5967 7098 5973 7100
rect 5727 7046 5729 7098
rect 5909 7046 5911 7098
rect 5665 7044 5671 7046
rect 5727 7044 5751 7046
rect 5807 7044 5831 7046
rect 5887 7044 5911 7046
rect 5967 7044 5973 7046
rect 5665 7035 5973 7044
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5828 6458 5856 6666
rect 6325 6556 6633 6565
rect 6325 6554 6331 6556
rect 6387 6554 6411 6556
rect 6467 6554 6491 6556
rect 6547 6554 6571 6556
rect 6627 6554 6633 6556
rect 6387 6502 6389 6554
rect 6569 6502 6571 6554
rect 6325 6500 6331 6502
rect 6387 6500 6411 6502
rect 6467 6500 6491 6502
rect 6547 6500 6571 6502
rect 6627 6500 6633 6502
rect 6325 6491 6633 6500
rect 6840 6458 6868 7346
rect 7551 7100 7859 7109
rect 7551 7098 7557 7100
rect 7613 7098 7637 7100
rect 7693 7098 7717 7100
rect 7773 7098 7797 7100
rect 7853 7098 7859 7100
rect 7613 7046 7615 7098
rect 7795 7046 7797 7098
rect 7551 7044 7557 7046
rect 7613 7044 7637 7046
rect 7693 7044 7717 7046
rect 7773 7044 7797 7046
rect 7853 7044 7859 7046
rect 7551 7035 7859 7044
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5552 5642 5580 6326
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 5665 6012 5973 6021
rect 5665 6010 5671 6012
rect 5727 6010 5751 6012
rect 5807 6010 5831 6012
rect 5887 6010 5911 6012
rect 5967 6010 5973 6012
rect 5727 5958 5729 6010
rect 5909 5958 5911 6010
rect 5665 5956 5671 5958
rect 5727 5956 5751 5958
rect 5807 5956 5831 5958
rect 5887 5956 5911 5958
rect 5967 5956 5973 5958
rect 5665 5947 5973 5956
rect 6012 5914 6040 6258
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6104 5794 6132 6190
rect 6012 5766 6132 5794
rect 6012 5642 6040 5766
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 6012 5370 6040 5578
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5908 5160 5960 5166
rect 6012 5114 6040 5306
rect 6196 5234 6224 6258
rect 7116 6186 7144 6598
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 7116 5574 7144 6122
rect 7551 6012 7859 6021
rect 7551 6010 7557 6012
rect 7613 6010 7637 6012
rect 7693 6010 7717 6012
rect 7773 6010 7797 6012
rect 7853 6010 7859 6012
rect 7613 5958 7615 6010
rect 7795 5958 7797 6010
rect 7551 5956 7557 5958
rect 7613 5956 7637 5958
rect 7693 5956 7717 5958
rect 7773 5956 7797 5958
rect 7853 5956 7859 5958
rect 7551 5947 7859 5956
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6325 5468 6633 5477
rect 6325 5466 6331 5468
rect 6387 5466 6411 5468
rect 6467 5466 6491 5468
rect 6547 5466 6571 5468
rect 6627 5466 6633 5468
rect 6387 5414 6389 5466
rect 6569 5414 6571 5466
rect 6325 5412 6331 5414
rect 6387 5412 6411 5414
rect 6467 5412 6491 5414
rect 6547 5412 6571 5414
rect 6627 5412 6633 5414
rect 6325 5403 6633 5412
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 5960 5108 6040 5114
rect 5908 5102 6040 5108
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 5920 5086 6040 5102
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4826 5580 4966
rect 5665 4924 5973 4933
rect 5665 4922 5671 4924
rect 5727 4922 5751 4924
rect 5807 4922 5831 4924
rect 5887 4922 5911 4924
rect 5967 4922 5973 4924
rect 5727 4870 5729 4922
rect 5909 4870 5911 4922
rect 5665 4868 5671 4870
rect 5727 4868 5751 4870
rect 5807 4868 5831 4870
rect 5887 4868 5911 4870
rect 5967 4868 5973 4870
rect 5665 4859 5973 4868
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 6012 4690 6040 5086
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6472 4554 6500 5102
rect 6656 4826 6684 5170
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4214 3280 4422
rect 4439 4380 4747 4389
rect 4439 4378 4445 4380
rect 4501 4378 4525 4380
rect 4581 4378 4605 4380
rect 4661 4378 4685 4380
rect 4741 4378 4747 4380
rect 4501 4326 4503 4378
rect 4683 4326 4685 4378
rect 4439 4324 4445 4326
rect 4501 4324 4525 4326
rect 4581 4324 4605 4326
rect 4661 4324 4685 4326
rect 4741 4324 4747 4326
rect 4439 4315 4747 4324
rect 6325 4380 6633 4389
rect 6325 4378 6331 4380
rect 6387 4378 6411 4380
rect 6467 4378 6491 4380
rect 6547 4378 6571 4380
rect 6627 4378 6633 4380
rect 6387 4326 6389 4378
rect 6569 4326 6571 4378
rect 6325 4324 6331 4326
rect 6387 4324 6411 4326
rect 6467 4324 6491 4326
rect 6547 4324 6571 4326
rect 6627 4324 6633 4326
rect 6325 4315 6633 4324
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 3779 3836 4087 3845
rect 3779 3834 3785 3836
rect 3841 3834 3865 3836
rect 3921 3834 3945 3836
rect 4001 3834 4025 3836
rect 4081 3834 4087 3836
rect 3841 3782 3843 3834
rect 4023 3782 4025 3834
rect 3779 3780 3785 3782
rect 3841 3780 3865 3782
rect 3921 3780 3945 3782
rect 4001 3780 4025 3782
rect 4081 3780 4087 3782
rect 3779 3771 4087 3780
rect 3779 2748 4087 2757
rect 3779 2746 3785 2748
rect 3841 2746 3865 2748
rect 3921 2746 3945 2748
rect 4001 2746 4025 2748
rect 4081 2746 4087 2748
rect 3841 2694 3843 2746
rect 4023 2694 4025 2746
rect 3779 2692 3785 2694
rect 3841 2692 3865 2694
rect 3921 2692 3945 2694
rect 4001 2692 4025 2694
rect 4081 2692 4087 2694
rect 3779 2683 4087 2692
rect 4264 2446 4292 3878
rect 5665 3836 5973 3845
rect 5665 3834 5671 3836
rect 5727 3834 5751 3836
rect 5807 3834 5831 3836
rect 5887 3834 5911 3836
rect 5967 3834 5973 3836
rect 5727 3782 5729 3834
rect 5909 3782 5911 3834
rect 5665 3780 5671 3782
rect 5727 3780 5751 3782
rect 5807 3780 5831 3782
rect 5887 3780 5911 3782
rect 5967 3780 5973 3782
rect 5665 3771 5973 3780
rect 4439 3292 4747 3301
rect 4439 3290 4445 3292
rect 4501 3290 4525 3292
rect 4581 3290 4605 3292
rect 4661 3290 4685 3292
rect 4741 3290 4747 3292
rect 4501 3238 4503 3290
rect 4683 3238 4685 3290
rect 4439 3236 4445 3238
rect 4501 3236 4525 3238
rect 4581 3236 4605 3238
rect 4661 3236 4685 3238
rect 4741 3236 4747 3238
rect 4439 3227 4747 3236
rect 6325 3292 6633 3301
rect 6325 3290 6331 3292
rect 6387 3290 6411 3292
rect 6467 3290 6491 3292
rect 6547 3290 6571 3292
rect 6627 3290 6633 3292
rect 6387 3238 6389 3290
rect 6569 3238 6571 3290
rect 6325 3236 6331 3238
rect 6387 3236 6411 3238
rect 6467 3236 6491 3238
rect 6547 3236 6571 3238
rect 6627 3236 6633 3238
rect 6325 3227 6633 3236
rect 6748 3126 6776 4558
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 5665 2748 5973 2757
rect 5665 2746 5671 2748
rect 5727 2746 5751 2748
rect 5807 2746 5831 2748
rect 5887 2746 5911 2748
rect 5967 2746 5973 2748
rect 5727 2694 5729 2746
rect 5909 2694 5911 2746
rect 5665 2692 5671 2694
rect 5727 2692 5751 2694
rect 5807 2692 5831 2694
rect 5887 2692 5911 2694
rect 5967 2692 5973 2694
rect 5665 2683 5973 2692
rect 7116 2446 7144 5510
rect 8128 5370 8156 8910
rect 8211 8732 8519 8741
rect 8211 8730 8217 8732
rect 8273 8730 8297 8732
rect 8353 8730 8377 8732
rect 8433 8730 8457 8732
rect 8513 8730 8519 8732
rect 8273 8678 8275 8730
rect 8455 8678 8457 8730
rect 8211 8676 8217 8678
rect 8273 8676 8297 8678
rect 8353 8676 8377 8678
rect 8433 8676 8457 8678
rect 8513 8676 8519 8678
rect 8211 8667 8519 8676
rect 8211 7644 8519 7653
rect 8211 7642 8217 7644
rect 8273 7642 8297 7644
rect 8353 7642 8377 7644
rect 8433 7642 8457 7644
rect 8513 7642 8519 7644
rect 8273 7590 8275 7642
rect 8455 7590 8457 7642
rect 8211 7588 8217 7590
rect 8273 7588 8297 7590
rect 8353 7588 8377 7590
rect 8433 7588 8457 7590
rect 8513 7588 8519 7590
rect 8211 7579 8519 7588
rect 8211 6556 8519 6565
rect 8211 6554 8217 6556
rect 8273 6554 8297 6556
rect 8353 6554 8377 6556
rect 8433 6554 8457 6556
rect 8513 6554 8519 6556
rect 8273 6502 8275 6554
rect 8455 6502 8457 6554
rect 8211 6500 8217 6502
rect 8273 6500 8297 6502
rect 8353 6500 8377 6502
rect 8433 6500 8457 6502
rect 8513 6500 8519 6502
rect 8211 6491 8519 6500
rect 8211 5468 8519 5477
rect 8211 5466 8217 5468
rect 8273 5466 8297 5468
rect 8353 5466 8377 5468
rect 8433 5466 8457 5468
rect 8513 5466 8519 5468
rect 8273 5414 8275 5466
rect 8455 5414 8457 5466
rect 8211 5412 8217 5414
rect 8273 5412 8297 5414
rect 8353 5412 8377 5414
rect 8433 5412 8457 5414
rect 8513 5412 8519 5414
rect 8211 5403 8519 5412
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7551 4924 7859 4933
rect 7551 4922 7557 4924
rect 7613 4922 7637 4924
rect 7693 4922 7717 4924
rect 7773 4922 7797 4924
rect 7853 4922 7859 4924
rect 7613 4870 7615 4922
rect 7795 4870 7797 4922
rect 7551 4868 7557 4870
rect 7613 4868 7637 4870
rect 7693 4868 7717 4870
rect 7773 4868 7797 4870
rect 7853 4868 7859 4870
rect 7551 4859 7859 4868
rect 8211 4380 8519 4389
rect 8211 4378 8217 4380
rect 8273 4378 8297 4380
rect 8353 4378 8377 4380
rect 8433 4378 8457 4380
rect 8513 4378 8519 4380
rect 8273 4326 8275 4378
rect 8455 4326 8457 4378
rect 8211 4324 8217 4326
rect 8273 4324 8297 4326
rect 8353 4324 8377 4326
rect 8433 4324 8457 4326
rect 8513 4324 8519 4326
rect 8211 4315 8519 4324
rect 7551 3836 7859 3845
rect 7551 3834 7557 3836
rect 7613 3834 7637 3836
rect 7693 3834 7717 3836
rect 7773 3834 7797 3836
rect 7853 3834 7859 3836
rect 7613 3782 7615 3834
rect 7795 3782 7797 3834
rect 7551 3780 7557 3782
rect 7613 3780 7637 3782
rect 7693 3780 7717 3782
rect 7773 3780 7797 3782
rect 7853 3780 7859 3782
rect 7551 3771 7859 3780
rect 8211 3292 8519 3301
rect 8211 3290 8217 3292
rect 8273 3290 8297 3292
rect 8353 3290 8377 3292
rect 8433 3290 8457 3292
rect 8513 3290 8519 3292
rect 8273 3238 8275 3290
rect 8455 3238 8457 3290
rect 8211 3236 8217 3238
rect 8273 3236 8297 3238
rect 8353 3236 8377 3238
rect 8433 3236 8457 3238
rect 8513 3236 8519 3238
rect 8211 3227 8519 3236
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8036 2825 8064 2994
rect 8022 2816 8078 2825
rect 7551 2748 7859 2757
rect 8022 2751 8078 2760
rect 7551 2746 7557 2748
rect 7613 2746 7637 2748
rect 7693 2746 7717 2748
rect 7773 2746 7797 2748
rect 7853 2746 7859 2748
rect 7613 2694 7615 2746
rect 7795 2694 7797 2746
rect 7551 2692 7557 2694
rect 7613 2692 7637 2694
rect 7693 2692 7717 2694
rect 7773 2692 7797 2694
rect 7853 2692 7859 2694
rect 7551 2683 7859 2692
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 32 800 60 2246
rect 2553 2204 2861 2213
rect 2553 2202 2559 2204
rect 2615 2202 2639 2204
rect 2695 2202 2719 2204
rect 2775 2202 2799 2204
rect 2855 2202 2861 2204
rect 2615 2150 2617 2202
rect 2797 2150 2799 2202
rect 2553 2148 2559 2150
rect 2615 2148 2639 2150
rect 2695 2148 2719 2150
rect 2775 2148 2799 2150
rect 2855 2148 2861 2150
rect 2553 2139 2861 2148
rect 3896 800 3924 2246
rect 4439 2204 4747 2213
rect 4439 2202 4445 2204
rect 4501 2202 4525 2204
rect 4581 2202 4605 2204
rect 4661 2202 4685 2204
rect 4741 2202 4747 2204
rect 4501 2150 4503 2202
rect 4683 2150 4685 2202
rect 4439 2148 4445 2150
rect 4501 2148 4525 2150
rect 4581 2148 4605 2150
rect 4661 2148 4685 2150
rect 4741 2148 4747 2150
rect 4439 2139 4747 2148
rect 6325 2204 6633 2213
rect 6325 2202 6331 2204
rect 6387 2202 6411 2204
rect 6467 2202 6491 2204
rect 6547 2202 6571 2204
rect 6627 2202 6633 2204
rect 6387 2150 6389 2202
rect 6569 2150 6571 2202
rect 6325 2148 6331 2150
rect 6387 2148 6411 2150
rect 6467 2148 6491 2150
rect 6547 2148 6571 2150
rect 6627 2148 6633 2150
rect 6325 2139 6633 2148
rect 8128 1442 8156 2246
rect 8211 2204 8519 2213
rect 8211 2202 8217 2204
rect 8273 2202 8297 2204
rect 8353 2202 8377 2204
rect 8433 2202 8457 2204
rect 8513 2202 8519 2204
rect 8273 2150 8275 2202
rect 8455 2150 8457 2202
rect 8211 2148 8217 2150
rect 8273 2148 8297 2150
rect 8353 2148 8377 2150
rect 8433 2148 8457 2150
rect 8513 2148 8519 2150
rect 8211 2139 8519 2148
rect 8128 1414 8432 1442
rect 8404 800 8432 1414
rect 18 0 74 800
rect 3882 0 3938 800
rect 8390 0 8446 800
<< via2 >>
rect 1899 9274 1955 9276
rect 1979 9274 2035 9276
rect 2059 9274 2115 9276
rect 2139 9274 2195 9276
rect 1899 9222 1945 9274
rect 1945 9222 1955 9274
rect 1979 9222 2009 9274
rect 2009 9222 2021 9274
rect 2021 9222 2035 9274
rect 2059 9222 2073 9274
rect 2073 9222 2085 9274
rect 2085 9222 2115 9274
rect 2139 9222 2149 9274
rect 2149 9222 2195 9274
rect 1899 9220 1955 9222
rect 1979 9220 2035 9222
rect 2059 9220 2115 9222
rect 2139 9220 2195 9222
rect 3785 9274 3841 9276
rect 3865 9274 3921 9276
rect 3945 9274 4001 9276
rect 4025 9274 4081 9276
rect 3785 9222 3831 9274
rect 3831 9222 3841 9274
rect 3865 9222 3895 9274
rect 3895 9222 3907 9274
rect 3907 9222 3921 9274
rect 3945 9222 3959 9274
rect 3959 9222 3971 9274
rect 3971 9222 4001 9274
rect 4025 9222 4035 9274
rect 4035 9222 4081 9274
rect 3785 9220 3841 9222
rect 3865 9220 3921 9222
rect 3945 9220 4001 9222
rect 4025 9220 4081 9222
rect 5671 9274 5727 9276
rect 5751 9274 5807 9276
rect 5831 9274 5887 9276
rect 5911 9274 5967 9276
rect 5671 9222 5717 9274
rect 5717 9222 5727 9274
rect 5751 9222 5781 9274
rect 5781 9222 5793 9274
rect 5793 9222 5807 9274
rect 5831 9222 5845 9274
rect 5845 9222 5857 9274
rect 5857 9222 5887 9274
rect 5911 9222 5921 9274
rect 5921 9222 5967 9274
rect 5671 9220 5727 9222
rect 5751 9220 5807 9222
rect 5831 9220 5887 9222
rect 5911 9220 5967 9222
rect 7557 9274 7613 9276
rect 7637 9274 7693 9276
rect 7717 9274 7773 9276
rect 7797 9274 7853 9276
rect 7557 9222 7603 9274
rect 7603 9222 7613 9274
rect 7637 9222 7667 9274
rect 7667 9222 7679 9274
rect 7679 9222 7693 9274
rect 7717 9222 7731 9274
rect 7731 9222 7743 9274
rect 7743 9222 7773 9274
rect 7797 9222 7807 9274
rect 7807 9222 7853 9274
rect 7557 9220 7613 9222
rect 7637 9220 7693 9222
rect 7717 9220 7773 9222
rect 7797 9220 7853 9222
rect 1766 8880 1822 8936
rect 2559 8730 2615 8732
rect 2639 8730 2695 8732
rect 2719 8730 2775 8732
rect 2799 8730 2855 8732
rect 2559 8678 2605 8730
rect 2605 8678 2615 8730
rect 2639 8678 2669 8730
rect 2669 8678 2681 8730
rect 2681 8678 2695 8730
rect 2719 8678 2733 8730
rect 2733 8678 2745 8730
rect 2745 8678 2775 8730
rect 2799 8678 2809 8730
rect 2809 8678 2855 8730
rect 2559 8676 2615 8678
rect 2639 8676 2695 8678
rect 2719 8676 2775 8678
rect 2799 8676 2855 8678
rect 4445 8730 4501 8732
rect 4525 8730 4581 8732
rect 4605 8730 4661 8732
rect 4685 8730 4741 8732
rect 4445 8678 4491 8730
rect 4491 8678 4501 8730
rect 4525 8678 4555 8730
rect 4555 8678 4567 8730
rect 4567 8678 4581 8730
rect 4605 8678 4619 8730
rect 4619 8678 4631 8730
rect 4631 8678 4661 8730
rect 4685 8678 4695 8730
rect 4695 8678 4741 8730
rect 4445 8676 4501 8678
rect 4525 8676 4581 8678
rect 4605 8676 4661 8678
rect 4685 8676 4741 8678
rect 1899 8186 1955 8188
rect 1979 8186 2035 8188
rect 2059 8186 2115 8188
rect 2139 8186 2195 8188
rect 1899 8134 1945 8186
rect 1945 8134 1955 8186
rect 1979 8134 2009 8186
rect 2009 8134 2021 8186
rect 2021 8134 2035 8186
rect 2059 8134 2073 8186
rect 2073 8134 2085 8186
rect 2085 8134 2115 8186
rect 2139 8134 2149 8186
rect 2149 8134 2195 8186
rect 1899 8132 1955 8134
rect 1979 8132 2035 8134
rect 2059 8132 2115 8134
rect 2139 8132 2195 8134
rect 3785 8186 3841 8188
rect 3865 8186 3921 8188
rect 3945 8186 4001 8188
rect 4025 8186 4081 8188
rect 3785 8134 3831 8186
rect 3831 8134 3841 8186
rect 3865 8134 3895 8186
rect 3895 8134 3907 8186
rect 3907 8134 3921 8186
rect 3945 8134 3959 8186
rect 3959 8134 3971 8186
rect 3971 8134 4001 8186
rect 4025 8134 4035 8186
rect 4035 8134 4081 8186
rect 3785 8132 3841 8134
rect 3865 8132 3921 8134
rect 3945 8132 4001 8134
rect 4025 8132 4081 8134
rect 2559 7642 2615 7644
rect 2639 7642 2695 7644
rect 2719 7642 2775 7644
rect 2799 7642 2855 7644
rect 2559 7590 2605 7642
rect 2605 7590 2615 7642
rect 2639 7590 2669 7642
rect 2669 7590 2681 7642
rect 2681 7590 2695 7642
rect 2719 7590 2733 7642
rect 2733 7590 2745 7642
rect 2745 7590 2775 7642
rect 2799 7590 2809 7642
rect 2809 7590 2855 7642
rect 2559 7588 2615 7590
rect 2639 7588 2695 7590
rect 2719 7588 2775 7590
rect 2799 7588 2855 7590
rect 1899 7098 1955 7100
rect 1979 7098 2035 7100
rect 2059 7098 2115 7100
rect 2139 7098 2195 7100
rect 1899 7046 1945 7098
rect 1945 7046 1955 7098
rect 1979 7046 2009 7098
rect 2009 7046 2021 7098
rect 2021 7046 2035 7098
rect 2059 7046 2073 7098
rect 2073 7046 2085 7098
rect 2085 7046 2115 7098
rect 2139 7046 2149 7098
rect 2149 7046 2195 7098
rect 1899 7044 1955 7046
rect 1979 7044 2035 7046
rect 2059 7044 2115 7046
rect 2139 7044 2195 7046
rect 3785 7098 3841 7100
rect 3865 7098 3921 7100
rect 3945 7098 4001 7100
rect 4025 7098 4081 7100
rect 3785 7046 3831 7098
rect 3831 7046 3841 7098
rect 3865 7046 3895 7098
rect 3895 7046 3907 7098
rect 3907 7046 3921 7098
rect 3945 7046 3959 7098
rect 3959 7046 3971 7098
rect 3971 7046 4001 7098
rect 4025 7046 4035 7098
rect 4035 7046 4081 7098
rect 3785 7044 3841 7046
rect 3865 7044 3921 7046
rect 3945 7044 4001 7046
rect 4025 7044 4081 7046
rect 2559 6554 2615 6556
rect 2639 6554 2695 6556
rect 2719 6554 2775 6556
rect 2799 6554 2855 6556
rect 2559 6502 2605 6554
rect 2605 6502 2615 6554
rect 2639 6502 2669 6554
rect 2669 6502 2681 6554
rect 2681 6502 2695 6554
rect 2719 6502 2733 6554
rect 2733 6502 2745 6554
rect 2745 6502 2775 6554
rect 2799 6502 2809 6554
rect 2809 6502 2855 6554
rect 2559 6500 2615 6502
rect 2639 6500 2695 6502
rect 2719 6500 2775 6502
rect 2799 6500 2855 6502
rect 1899 6010 1955 6012
rect 1979 6010 2035 6012
rect 2059 6010 2115 6012
rect 2139 6010 2195 6012
rect 1899 5958 1945 6010
rect 1945 5958 1955 6010
rect 1979 5958 2009 6010
rect 2009 5958 2021 6010
rect 2021 5958 2035 6010
rect 2059 5958 2073 6010
rect 2073 5958 2085 6010
rect 2085 5958 2115 6010
rect 2139 5958 2149 6010
rect 2149 5958 2195 6010
rect 1899 5956 1955 5958
rect 1979 5956 2035 5958
rect 2059 5956 2115 5958
rect 2139 5956 2195 5958
rect 3785 6010 3841 6012
rect 3865 6010 3921 6012
rect 3945 6010 4001 6012
rect 4025 6010 4081 6012
rect 3785 5958 3831 6010
rect 3831 5958 3841 6010
rect 3865 5958 3895 6010
rect 3895 5958 3907 6010
rect 3907 5958 3921 6010
rect 3945 5958 3959 6010
rect 3959 5958 3971 6010
rect 3971 5958 4001 6010
rect 4025 5958 4035 6010
rect 4035 5958 4081 6010
rect 3785 5956 3841 5958
rect 3865 5956 3921 5958
rect 3945 5956 4001 5958
rect 4025 5956 4081 5958
rect 4445 7642 4501 7644
rect 4525 7642 4581 7644
rect 4605 7642 4661 7644
rect 4685 7642 4741 7644
rect 4445 7590 4491 7642
rect 4491 7590 4501 7642
rect 4525 7590 4555 7642
rect 4555 7590 4567 7642
rect 4567 7590 4581 7642
rect 4605 7590 4619 7642
rect 4619 7590 4631 7642
rect 4631 7590 4661 7642
rect 4685 7590 4695 7642
rect 4695 7590 4741 7642
rect 4445 7588 4501 7590
rect 4525 7588 4581 7590
rect 4605 7588 4661 7590
rect 4685 7588 4741 7590
rect 4445 6554 4501 6556
rect 4525 6554 4581 6556
rect 4605 6554 4661 6556
rect 4685 6554 4741 6556
rect 4445 6502 4491 6554
rect 4491 6502 4501 6554
rect 4525 6502 4555 6554
rect 4555 6502 4567 6554
rect 4567 6502 4581 6554
rect 4605 6502 4619 6554
rect 4619 6502 4631 6554
rect 4631 6502 4661 6554
rect 4685 6502 4695 6554
rect 4695 6502 4741 6554
rect 4445 6500 4501 6502
rect 4525 6500 4581 6502
rect 4605 6500 4661 6502
rect 4685 6500 4741 6502
rect 2559 5466 2615 5468
rect 2639 5466 2695 5468
rect 2719 5466 2775 5468
rect 2799 5466 2855 5468
rect 2559 5414 2605 5466
rect 2605 5414 2615 5466
rect 2639 5414 2669 5466
rect 2669 5414 2681 5466
rect 2681 5414 2695 5466
rect 2719 5414 2733 5466
rect 2733 5414 2745 5466
rect 2745 5414 2775 5466
rect 2799 5414 2809 5466
rect 2809 5414 2855 5466
rect 2559 5412 2615 5414
rect 2639 5412 2695 5414
rect 2719 5412 2775 5414
rect 2799 5412 2855 5414
rect 4445 5466 4501 5468
rect 4525 5466 4581 5468
rect 4605 5466 4661 5468
rect 4685 5466 4741 5468
rect 4445 5414 4491 5466
rect 4491 5414 4501 5466
rect 4525 5414 4555 5466
rect 4555 5414 4567 5466
rect 4567 5414 4581 5466
rect 4605 5414 4619 5466
rect 4619 5414 4631 5466
rect 4631 5414 4661 5466
rect 4685 5414 4695 5466
rect 4695 5414 4741 5466
rect 4445 5412 4501 5414
rect 4525 5412 4581 5414
rect 4605 5412 4661 5414
rect 4685 5412 4741 5414
rect 6331 8730 6387 8732
rect 6411 8730 6467 8732
rect 6491 8730 6547 8732
rect 6571 8730 6627 8732
rect 6331 8678 6377 8730
rect 6377 8678 6387 8730
rect 6411 8678 6441 8730
rect 6441 8678 6453 8730
rect 6453 8678 6467 8730
rect 6491 8678 6505 8730
rect 6505 8678 6517 8730
rect 6517 8678 6547 8730
rect 6571 8678 6581 8730
rect 6581 8678 6627 8730
rect 6331 8676 6387 8678
rect 6411 8676 6467 8678
rect 6491 8676 6547 8678
rect 6571 8676 6627 8678
rect 5671 8186 5727 8188
rect 5751 8186 5807 8188
rect 5831 8186 5887 8188
rect 5911 8186 5967 8188
rect 5671 8134 5717 8186
rect 5717 8134 5727 8186
rect 5751 8134 5781 8186
rect 5781 8134 5793 8186
rect 5793 8134 5807 8186
rect 5831 8134 5845 8186
rect 5845 8134 5857 8186
rect 5857 8134 5887 8186
rect 5911 8134 5921 8186
rect 5921 8134 5967 8186
rect 5671 8132 5727 8134
rect 5751 8132 5807 8134
rect 5831 8132 5887 8134
rect 5911 8132 5967 8134
rect 7557 8186 7613 8188
rect 7637 8186 7693 8188
rect 7717 8186 7773 8188
rect 7797 8186 7853 8188
rect 7557 8134 7603 8186
rect 7603 8134 7613 8186
rect 7637 8134 7667 8186
rect 7667 8134 7679 8186
rect 7679 8134 7693 8186
rect 7717 8134 7731 8186
rect 7731 8134 7743 8186
rect 7743 8134 7773 8186
rect 7797 8134 7807 8186
rect 7807 8134 7853 8186
rect 7557 8132 7613 8134
rect 7637 8132 7693 8134
rect 7717 8132 7773 8134
rect 7797 8132 7853 8134
rect 6331 7642 6387 7644
rect 6411 7642 6467 7644
rect 6491 7642 6547 7644
rect 6571 7642 6627 7644
rect 6331 7590 6377 7642
rect 6377 7590 6387 7642
rect 6411 7590 6441 7642
rect 6441 7590 6453 7642
rect 6453 7590 6467 7642
rect 6491 7590 6505 7642
rect 6505 7590 6517 7642
rect 6517 7590 6547 7642
rect 6571 7590 6581 7642
rect 6581 7590 6627 7642
rect 6331 7588 6387 7590
rect 6411 7588 6467 7590
rect 6491 7588 6547 7590
rect 6571 7588 6627 7590
rect 1899 4922 1955 4924
rect 1979 4922 2035 4924
rect 2059 4922 2115 4924
rect 2139 4922 2195 4924
rect 1899 4870 1945 4922
rect 1945 4870 1955 4922
rect 1979 4870 2009 4922
rect 2009 4870 2021 4922
rect 2021 4870 2035 4922
rect 2059 4870 2073 4922
rect 2073 4870 2085 4922
rect 2085 4870 2115 4922
rect 2139 4870 2149 4922
rect 2149 4870 2195 4922
rect 1899 4868 1955 4870
rect 1979 4868 2035 4870
rect 2059 4868 2115 4870
rect 2139 4868 2195 4870
rect 2559 4378 2615 4380
rect 2639 4378 2695 4380
rect 2719 4378 2775 4380
rect 2799 4378 2855 4380
rect 2559 4326 2605 4378
rect 2605 4326 2615 4378
rect 2639 4326 2669 4378
rect 2669 4326 2681 4378
rect 2681 4326 2695 4378
rect 2719 4326 2733 4378
rect 2733 4326 2745 4378
rect 2745 4326 2775 4378
rect 2799 4326 2809 4378
rect 2809 4326 2855 4378
rect 2559 4324 2615 4326
rect 2639 4324 2695 4326
rect 2719 4324 2775 4326
rect 2799 4324 2855 4326
rect 1674 4120 1730 4176
rect 1899 3834 1955 3836
rect 1979 3834 2035 3836
rect 2059 3834 2115 3836
rect 2139 3834 2195 3836
rect 1899 3782 1945 3834
rect 1945 3782 1955 3834
rect 1979 3782 2009 3834
rect 2009 3782 2021 3834
rect 2021 3782 2035 3834
rect 2059 3782 2073 3834
rect 2073 3782 2085 3834
rect 2085 3782 2115 3834
rect 2139 3782 2149 3834
rect 2149 3782 2195 3834
rect 1899 3780 1955 3782
rect 1979 3780 2035 3782
rect 2059 3780 2115 3782
rect 2139 3780 2195 3782
rect 2559 3290 2615 3292
rect 2639 3290 2695 3292
rect 2719 3290 2775 3292
rect 2799 3290 2855 3292
rect 2559 3238 2605 3290
rect 2605 3238 2615 3290
rect 2639 3238 2669 3290
rect 2669 3238 2681 3290
rect 2681 3238 2695 3290
rect 2719 3238 2733 3290
rect 2733 3238 2745 3290
rect 2745 3238 2775 3290
rect 2799 3238 2809 3290
rect 2809 3238 2855 3290
rect 2559 3236 2615 3238
rect 2639 3236 2695 3238
rect 2719 3236 2775 3238
rect 2799 3236 2855 3238
rect 1899 2746 1955 2748
rect 1979 2746 2035 2748
rect 2059 2746 2115 2748
rect 2139 2746 2195 2748
rect 1899 2694 1945 2746
rect 1945 2694 1955 2746
rect 1979 2694 2009 2746
rect 2009 2694 2021 2746
rect 2021 2694 2035 2746
rect 2059 2694 2073 2746
rect 2073 2694 2085 2746
rect 2085 2694 2115 2746
rect 2139 2694 2149 2746
rect 2149 2694 2195 2746
rect 1899 2692 1955 2694
rect 1979 2692 2035 2694
rect 2059 2692 2115 2694
rect 2139 2692 2195 2694
rect 3785 4922 3841 4924
rect 3865 4922 3921 4924
rect 3945 4922 4001 4924
rect 4025 4922 4081 4924
rect 3785 4870 3831 4922
rect 3831 4870 3841 4922
rect 3865 4870 3895 4922
rect 3895 4870 3907 4922
rect 3907 4870 3921 4922
rect 3945 4870 3959 4922
rect 3959 4870 3971 4922
rect 3971 4870 4001 4922
rect 4025 4870 4035 4922
rect 4035 4870 4081 4922
rect 3785 4868 3841 4870
rect 3865 4868 3921 4870
rect 3945 4868 4001 4870
rect 4025 4868 4081 4870
rect 8022 7384 8078 7440
rect 5671 7098 5727 7100
rect 5751 7098 5807 7100
rect 5831 7098 5887 7100
rect 5911 7098 5967 7100
rect 5671 7046 5717 7098
rect 5717 7046 5727 7098
rect 5751 7046 5781 7098
rect 5781 7046 5793 7098
rect 5793 7046 5807 7098
rect 5831 7046 5845 7098
rect 5845 7046 5857 7098
rect 5857 7046 5887 7098
rect 5911 7046 5921 7098
rect 5921 7046 5967 7098
rect 5671 7044 5727 7046
rect 5751 7044 5807 7046
rect 5831 7044 5887 7046
rect 5911 7044 5967 7046
rect 6331 6554 6387 6556
rect 6411 6554 6467 6556
rect 6491 6554 6547 6556
rect 6571 6554 6627 6556
rect 6331 6502 6377 6554
rect 6377 6502 6387 6554
rect 6411 6502 6441 6554
rect 6441 6502 6453 6554
rect 6453 6502 6467 6554
rect 6491 6502 6505 6554
rect 6505 6502 6517 6554
rect 6517 6502 6547 6554
rect 6571 6502 6581 6554
rect 6581 6502 6627 6554
rect 6331 6500 6387 6502
rect 6411 6500 6467 6502
rect 6491 6500 6547 6502
rect 6571 6500 6627 6502
rect 7557 7098 7613 7100
rect 7637 7098 7693 7100
rect 7717 7098 7773 7100
rect 7797 7098 7853 7100
rect 7557 7046 7603 7098
rect 7603 7046 7613 7098
rect 7637 7046 7667 7098
rect 7667 7046 7679 7098
rect 7679 7046 7693 7098
rect 7717 7046 7731 7098
rect 7731 7046 7743 7098
rect 7743 7046 7773 7098
rect 7797 7046 7807 7098
rect 7807 7046 7853 7098
rect 7557 7044 7613 7046
rect 7637 7044 7693 7046
rect 7717 7044 7773 7046
rect 7797 7044 7853 7046
rect 5671 6010 5727 6012
rect 5751 6010 5807 6012
rect 5831 6010 5887 6012
rect 5911 6010 5967 6012
rect 5671 5958 5717 6010
rect 5717 5958 5727 6010
rect 5751 5958 5781 6010
rect 5781 5958 5793 6010
rect 5793 5958 5807 6010
rect 5831 5958 5845 6010
rect 5845 5958 5857 6010
rect 5857 5958 5887 6010
rect 5911 5958 5921 6010
rect 5921 5958 5967 6010
rect 5671 5956 5727 5958
rect 5751 5956 5807 5958
rect 5831 5956 5887 5958
rect 5911 5956 5967 5958
rect 7557 6010 7613 6012
rect 7637 6010 7693 6012
rect 7717 6010 7773 6012
rect 7797 6010 7853 6012
rect 7557 5958 7603 6010
rect 7603 5958 7613 6010
rect 7637 5958 7667 6010
rect 7667 5958 7679 6010
rect 7679 5958 7693 6010
rect 7717 5958 7731 6010
rect 7731 5958 7743 6010
rect 7743 5958 7773 6010
rect 7797 5958 7807 6010
rect 7807 5958 7853 6010
rect 7557 5956 7613 5958
rect 7637 5956 7693 5958
rect 7717 5956 7773 5958
rect 7797 5956 7853 5958
rect 6331 5466 6387 5468
rect 6411 5466 6467 5468
rect 6491 5466 6547 5468
rect 6571 5466 6627 5468
rect 6331 5414 6377 5466
rect 6377 5414 6387 5466
rect 6411 5414 6441 5466
rect 6441 5414 6453 5466
rect 6453 5414 6467 5466
rect 6491 5414 6505 5466
rect 6505 5414 6517 5466
rect 6517 5414 6547 5466
rect 6571 5414 6581 5466
rect 6581 5414 6627 5466
rect 6331 5412 6387 5414
rect 6411 5412 6467 5414
rect 6491 5412 6547 5414
rect 6571 5412 6627 5414
rect 5671 4922 5727 4924
rect 5751 4922 5807 4924
rect 5831 4922 5887 4924
rect 5911 4922 5967 4924
rect 5671 4870 5717 4922
rect 5717 4870 5727 4922
rect 5751 4870 5781 4922
rect 5781 4870 5793 4922
rect 5793 4870 5807 4922
rect 5831 4870 5845 4922
rect 5845 4870 5857 4922
rect 5857 4870 5887 4922
rect 5911 4870 5921 4922
rect 5921 4870 5967 4922
rect 5671 4868 5727 4870
rect 5751 4868 5807 4870
rect 5831 4868 5887 4870
rect 5911 4868 5967 4870
rect 4445 4378 4501 4380
rect 4525 4378 4581 4380
rect 4605 4378 4661 4380
rect 4685 4378 4741 4380
rect 4445 4326 4491 4378
rect 4491 4326 4501 4378
rect 4525 4326 4555 4378
rect 4555 4326 4567 4378
rect 4567 4326 4581 4378
rect 4605 4326 4619 4378
rect 4619 4326 4631 4378
rect 4631 4326 4661 4378
rect 4685 4326 4695 4378
rect 4695 4326 4741 4378
rect 4445 4324 4501 4326
rect 4525 4324 4581 4326
rect 4605 4324 4661 4326
rect 4685 4324 4741 4326
rect 6331 4378 6387 4380
rect 6411 4378 6467 4380
rect 6491 4378 6547 4380
rect 6571 4378 6627 4380
rect 6331 4326 6377 4378
rect 6377 4326 6387 4378
rect 6411 4326 6441 4378
rect 6441 4326 6453 4378
rect 6453 4326 6467 4378
rect 6491 4326 6505 4378
rect 6505 4326 6517 4378
rect 6517 4326 6547 4378
rect 6571 4326 6581 4378
rect 6581 4326 6627 4378
rect 6331 4324 6387 4326
rect 6411 4324 6467 4326
rect 6491 4324 6547 4326
rect 6571 4324 6627 4326
rect 3785 3834 3841 3836
rect 3865 3834 3921 3836
rect 3945 3834 4001 3836
rect 4025 3834 4081 3836
rect 3785 3782 3831 3834
rect 3831 3782 3841 3834
rect 3865 3782 3895 3834
rect 3895 3782 3907 3834
rect 3907 3782 3921 3834
rect 3945 3782 3959 3834
rect 3959 3782 3971 3834
rect 3971 3782 4001 3834
rect 4025 3782 4035 3834
rect 4035 3782 4081 3834
rect 3785 3780 3841 3782
rect 3865 3780 3921 3782
rect 3945 3780 4001 3782
rect 4025 3780 4081 3782
rect 3785 2746 3841 2748
rect 3865 2746 3921 2748
rect 3945 2746 4001 2748
rect 4025 2746 4081 2748
rect 3785 2694 3831 2746
rect 3831 2694 3841 2746
rect 3865 2694 3895 2746
rect 3895 2694 3907 2746
rect 3907 2694 3921 2746
rect 3945 2694 3959 2746
rect 3959 2694 3971 2746
rect 3971 2694 4001 2746
rect 4025 2694 4035 2746
rect 4035 2694 4081 2746
rect 3785 2692 3841 2694
rect 3865 2692 3921 2694
rect 3945 2692 4001 2694
rect 4025 2692 4081 2694
rect 5671 3834 5727 3836
rect 5751 3834 5807 3836
rect 5831 3834 5887 3836
rect 5911 3834 5967 3836
rect 5671 3782 5717 3834
rect 5717 3782 5727 3834
rect 5751 3782 5781 3834
rect 5781 3782 5793 3834
rect 5793 3782 5807 3834
rect 5831 3782 5845 3834
rect 5845 3782 5857 3834
rect 5857 3782 5887 3834
rect 5911 3782 5921 3834
rect 5921 3782 5967 3834
rect 5671 3780 5727 3782
rect 5751 3780 5807 3782
rect 5831 3780 5887 3782
rect 5911 3780 5967 3782
rect 4445 3290 4501 3292
rect 4525 3290 4581 3292
rect 4605 3290 4661 3292
rect 4685 3290 4741 3292
rect 4445 3238 4491 3290
rect 4491 3238 4501 3290
rect 4525 3238 4555 3290
rect 4555 3238 4567 3290
rect 4567 3238 4581 3290
rect 4605 3238 4619 3290
rect 4619 3238 4631 3290
rect 4631 3238 4661 3290
rect 4685 3238 4695 3290
rect 4695 3238 4741 3290
rect 4445 3236 4501 3238
rect 4525 3236 4581 3238
rect 4605 3236 4661 3238
rect 4685 3236 4741 3238
rect 6331 3290 6387 3292
rect 6411 3290 6467 3292
rect 6491 3290 6547 3292
rect 6571 3290 6627 3292
rect 6331 3238 6377 3290
rect 6377 3238 6387 3290
rect 6411 3238 6441 3290
rect 6441 3238 6453 3290
rect 6453 3238 6467 3290
rect 6491 3238 6505 3290
rect 6505 3238 6517 3290
rect 6517 3238 6547 3290
rect 6571 3238 6581 3290
rect 6581 3238 6627 3290
rect 6331 3236 6387 3238
rect 6411 3236 6467 3238
rect 6491 3236 6547 3238
rect 6571 3236 6627 3238
rect 5671 2746 5727 2748
rect 5751 2746 5807 2748
rect 5831 2746 5887 2748
rect 5911 2746 5967 2748
rect 5671 2694 5717 2746
rect 5717 2694 5727 2746
rect 5751 2694 5781 2746
rect 5781 2694 5793 2746
rect 5793 2694 5807 2746
rect 5831 2694 5845 2746
rect 5845 2694 5857 2746
rect 5857 2694 5887 2746
rect 5911 2694 5921 2746
rect 5921 2694 5967 2746
rect 5671 2692 5727 2694
rect 5751 2692 5807 2694
rect 5831 2692 5887 2694
rect 5911 2692 5967 2694
rect 8217 8730 8273 8732
rect 8297 8730 8353 8732
rect 8377 8730 8433 8732
rect 8457 8730 8513 8732
rect 8217 8678 8263 8730
rect 8263 8678 8273 8730
rect 8297 8678 8327 8730
rect 8327 8678 8339 8730
rect 8339 8678 8353 8730
rect 8377 8678 8391 8730
rect 8391 8678 8403 8730
rect 8403 8678 8433 8730
rect 8457 8678 8467 8730
rect 8467 8678 8513 8730
rect 8217 8676 8273 8678
rect 8297 8676 8353 8678
rect 8377 8676 8433 8678
rect 8457 8676 8513 8678
rect 8217 7642 8273 7644
rect 8297 7642 8353 7644
rect 8377 7642 8433 7644
rect 8457 7642 8513 7644
rect 8217 7590 8263 7642
rect 8263 7590 8273 7642
rect 8297 7590 8327 7642
rect 8327 7590 8339 7642
rect 8339 7590 8353 7642
rect 8377 7590 8391 7642
rect 8391 7590 8403 7642
rect 8403 7590 8433 7642
rect 8457 7590 8467 7642
rect 8467 7590 8513 7642
rect 8217 7588 8273 7590
rect 8297 7588 8353 7590
rect 8377 7588 8433 7590
rect 8457 7588 8513 7590
rect 8217 6554 8273 6556
rect 8297 6554 8353 6556
rect 8377 6554 8433 6556
rect 8457 6554 8513 6556
rect 8217 6502 8263 6554
rect 8263 6502 8273 6554
rect 8297 6502 8327 6554
rect 8327 6502 8339 6554
rect 8339 6502 8353 6554
rect 8377 6502 8391 6554
rect 8391 6502 8403 6554
rect 8403 6502 8433 6554
rect 8457 6502 8467 6554
rect 8467 6502 8513 6554
rect 8217 6500 8273 6502
rect 8297 6500 8353 6502
rect 8377 6500 8433 6502
rect 8457 6500 8513 6502
rect 8217 5466 8273 5468
rect 8297 5466 8353 5468
rect 8377 5466 8433 5468
rect 8457 5466 8513 5468
rect 8217 5414 8263 5466
rect 8263 5414 8273 5466
rect 8297 5414 8327 5466
rect 8327 5414 8339 5466
rect 8339 5414 8353 5466
rect 8377 5414 8391 5466
rect 8391 5414 8403 5466
rect 8403 5414 8433 5466
rect 8457 5414 8467 5466
rect 8467 5414 8513 5466
rect 8217 5412 8273 5414
rect 8297 5412 8353 5414
rect 8377 5412 8433 5414
rect 8457 5412 8513 5414
rect 7557 4922 7613 4924
rect 7637 4922 7693 4924
rect 7717 4922 7773 4924
rect 7797 4922 7853 4924
rect 7557 4870 7603 4922
rect 7603 4870 7613 4922
rect 7637 4870 7667 4922
rect 7667 4870 7679 4922
rect 7679 4870 7693 4922
rect 7717 4870 7731 4922
rect 7731 4870 7743 4922
rect 7743 4870 7773 4922
rect 7797 4870 7807 4922
rect 7807 4870 7853 4922
rect 7557 4868 7613 4870
rect 7637 4868 7693 4870
rect 7717 4868 7773 4870
rect 7797 4868 7853 4870
rect 8217 4378 8273 4380
rect 8297 4378 8353 4380
rect 8377 4378 8433 4380
rect 8457 4378 8513 4380
rect 8217 4326 8263 4378
rect 8263 4326 8273 4378
rect 8297 4326 8327 4378
rect 8327 4326 8339 4378
rect 8339 4326 8353 4378
rect 8377 4326 8391 4378
rect 8391 4326 8403 4378
rect 8403 4326 8433 4378
rect 8457 4326 8467 4378
rect 8467 4326 8513 4378
rect 8217 4324 8273 4326
rect 8297 4324 8353 4326
rect 8377 4324 8433 4326
rect 8457 4324 8513 4326
rect 7557 3834 7613 3836
rect 7637 3834 7693 3836
rect 7717 3834 7773 3836
rect 7797 3834 7853 3836
rect 7557 3782 7603 3834
rect 7603 3782 7613 3834
rect 7637 3782 7667 3834
rect 7667 3782 7679 3834
rect 7679 3782 7693 3834
rect 7717 3782 7731 3834
rect 7731 3782 7743 3834
rect 7743 3782 7773 3834
rect 7797 3782 7807 3834
rect 7807 3782 7853 3834
rect 7557 3780 7613 3782
rect 7637 3780 7693 3782
rect 7717 3780 7773 3782
rect 7797 3780 7853 3782
rect 8217 3290 8273 3292
rect 8297 3290 8353 3292
rect 8377 3290 8433 3292
rect 8457 3290 8513 3292
rect 8217 3238 8263 3290
rect 8263 3238 8273 3290
rect 8297 3238 8327 3290
rect 8327 3238 8339 3290
rect 8339 3238 8353 3290
rect 8377 3238 8391 3290
rect 8391 3238 8403 3290
rect 8403 3238 8433 3290
rect 8457 3238 8467 3290
rect 8467 3238 8513 3290
rect 8217 3236 8273 3238
rect 8297 3236 8353 3238
rect 8377 3236 8433 3238
rect 8457 3236 8513 3238
rect 8022 2760 8078 2816
rect 7557 2746 7613 2748
rect 7637 2746 7693 2748
rect 7717 2746 7773 2748
rect 7797 2746 7853 2748
rect 7557 2694 7603 2746
rect 7603 2694 7613 2746
rect 7637 2694 7667 2746
rect 7667 2694 7679 2746
rect 7679 2694 7693 2746
rect 7717 2694 7731 2746
rect 7731 2694 7743 2746
rect 7743 2694 7773 2746
rect 7797 2694 7807 2746
rect 7807 2694 7853 2746
rect 7557 2692 7613 2694
rect 7637 2692 7693 2694
rect 7717 2692 7773 2694
rect 7797 2692 7853 2694
rect 2559 2202 2615 2204
rect 2639 2202 2695 2204
rect 2719 2202 2775 2204
rect 2799 2202 2855 2204
rect 2559 2150 2605 2202
rect 2605 2150 2615 2202
rect 2639 2150 2669 2202
rect 2669 2150 2681 2202
rect 2681 2150 2695 2202
rect 2719 2150 2733 2202
rect 2733 2150 2745 2202
rect 2745 2150 2775 2202
rect 2799 2150 2809 2202
rect 2809 2150 2855 2202
rect 2559 2148 2615 2150
rect 2639 2148 2695 2150
rect 2719 2148 2775 2150
rect 2799 2148 2855 2150
rect 4445 2202 4501 2204
rect 4525 2202 4581 2204
rect 4605 2202 4661 2204
rect 4685 2202 4741 2204
rect 4445 2150 4491 2202
rect 4491 2150 4501 2202
rect 4525 2150 4555 2202
rect 4555 2150 4567 2202
rect 4567 2150 4581 2202
rect 4605 2150 4619 2202
rect 4619 2150 4631 2202
rect 4631 2150 4661 2202
rect 4685 2150 4695 2202
rect 4695 2150 4741 2202
rect 4445 2148 4501 2150
rect 4525 2148 4581 2150
rect 4605 2148 4661 2150
rect 4685 2148 4741 2150
rect 6331 2202 6387 2204
rect 6411 2202 6467 2204
rect 6491 2202 6547 2204
rect 6571 2202 6627 2204
rect 6331 2150 6377 2202
rect 6377 2150 6387 2202
rect 6411 2150 6441 2202
rect 6441 2150 6453 2202
rect 6453 2150 6467 2202
rect 6491 2150 6505 2202
rect 6505 2150 6517 2202
rect 6517 2150 6547 2202
rect 6571 2150 6581 2202
rect 6581 2150 6627 2202
rect 6331 2148 6387 2150
rect 6411 2148 6467 2150
rect 6491 2148 6547 2150
rect 6571 2148 6627 2150
rect 8217 2202 8273 2204
rect 8297 2202 8353 2204
rect 8377 2202 8433 2204
rect 8457 2202 8513 2204
rect 8217 2150 8263 2202
rect 8263 2150 8273 2202
rect 8297 2150 8327 2202
rect 8327 2150 8339 2202
rect 8339 2150 8353 2202
rect 8377 2150 8391 2202
rect 8391 2150 8403 2202
rect 8403 2150 8433 2202
rect 8457 2150 8467 2202
rect 8467 2150 8513 2202
rect 8217 2148 8273 2150
rect 8297 2148 8353 2150
rect 8377 2148 8433 2150
rect 8457 2148 8513 2150
<< metal3 >>
rect 1889 9280 2205 9281
rect 1889 9216 1895 9280
rect 1959 9216 1975 9280
rect 2039 9216 2055 9280
rect 2119 9216 2135 9280
rect 2199 9216 2205 9280
rect 1889 9215 2205 9216
rect 3775 9280 4091 9281
rect 3775 9216 3781 9280
rect 3845 9216 3861 9280
rect 3925 9216 3941 9280
rect 4005 9216 4021 9280
rect 4085 9216 4091 9280
rect 3775 9215 4091 9216
rect 5661 9280 5977 9281
rect 5661 9216 5667 9280
rect 5731 9216 5747 9280
rect 5811 9216 5827 9280
rect 5891 9216 5907 9280
rect 5971 9216 5977 9280
rect 5661 9215 5977 9216
rect 7547 9280 7863 9281
rect 7547 9216 7553 9280
rect 7617 9216 7633 9280
rect 7697 9216 7713 9280
rect 7777 9216 7793 9280
rect 7857 9216 7863 9280
rect 7547 9215 7863 9216
rect 0 8938 800 8968
rect 1761 8938 1827 8941
rect 0 8936 1827 8938
rect 0 8880 1766 8936
rect 1822 8880 1827 8936
rect 0 8878 1827 8880
rect 0 8848 800 8878
rect 1761 8875 1827 8878
rect 2549 8736 2865 8737
rect 2549 8672 2555 8736
rect 2619 8672 2635 8736
rect 2699 8672 2715 8736
rect 2779 8672 2795 8736
rect 2859 8672 2865 8736
rect 2549 8671 2865 8672
rect 4435 8736 4751 8737
rect 4435 8672 4441 8736
rect 4505 8672 4521 8736
rect 4585 8672 4601 8736
rect 4665 8672 4681 8736
rect 4745 8672 4751 8736
rect 4435 8671 4751 8672
rect 6321 8736 6637 8737
rect 6321 8672 6327 8736
rect 6391 8672 6407 8736
rect 6471 8672 6487 8736
rect 6551 8672 6567 8736
rect 6631 8672 6637 8736
rect 6321 8671 6637 8672
rect 8207 8736 8523 8737
rect 8207 8672 8213 8736
rect 8277 8672 8293 8736
rect 8357 8672 8373 8736
rect 8437 8672 8453 8736
rect 8517 8672 8523 8736
rect 8207 8671 8523 8672
rect 1889 8192 2205 8193
rect 1889 8128 1895 8192
rect 1959 8128 1975 8192
rect 2039 8128 2055 8192
rect 2119 8128 2135 8192
rect 2199 8128 2205 8192
rect 1889 8127 2205 8128
rect 3775 8192 4091 8193
rect 3775 8128 3781 8192
rect 3845 8128 3861 8192
rect 3925 8128 3941 8192
rect 4005 8128 4021 8192
rect 4085 8128 4091 8192
rect 3775 8127 4091 8128
rect 5661 8192 5977 8193
rect 5661 8128 5667 8192
rect 5731 8128 5747 8192
rect 5811 8128 5827 8192
rect 5891 8128 5907 8192
rect 5971 8128 5977 8192
rect 5661 8127 5977 8128
rect 7547 8192 7863 8193
rect 7547 8128 7553 8192
rect 7617 8128 7633 8192
rect 7697 8128 7713 8192
rect 7777 8128 7793 8192
rect 7857 8128 7863 8192
rect 7547 8127 7863 8128
rect 2549 7648 2865 7649
rect 2549 7584 2555 7648
rect 2619 7584 2635 7648
rect 2699 7584 2715 7648
rect 2779 7584 2795 7648
rect 2859 7584 2865 7648
rect 2549 7583 2865 7584
rect 4435 7648 4751 7649
rect 4435 7584 4441 7648
rect 4505 7584 4521 7648
rect 4585 7584 4601 7648
rect 4665 7584 4681 7648
rect 4745 7584 4751 7648
rect 4435 7583 4751 7584
rect 6321 7648 6637 7649
rect 6321 7584 6327 7648
rect 6391 7584 6407 7648
rect 6471 7584 6487 7648
rect 6551 7584 6567 7648
rect 6631 7584 6637 7648
rect 6321 7583 6637 7584
rect 8207 7648 8523 7649
rect 8207 7584 8213 7648
rect 8277 7584 8293 7648
rect 8357 7584 8373 7648
rect 8437 7584 8453 7648
rect 8517 7584 8523 7648
rect 8207 7583 8523 7584
rect 8978 7578 9778 7608
rect 8710 7518 9778 7578
rect 8017 7442 8083 7445
rect 8710 7442 8770 7518
rect 8978 7488 9778 7518
rect 8017 7440 8770 7442
rect 8017 7384 8022 7440
rect 8078 7384 8770 7440
rect 8017 7382 8770 7384
rect 8017 7379 8083 7382
rect 1889 7104 2205 7105
rect 1889 7040 1895 7104
rect 1959 7040 1975 7104
rect 2039 7040 2055 7104
rect 2119 7040 2135 7104
rect 2199 7040 2205 7104
rect 1889 7039 2205 7040
rect 3775 7104 4091 7105
rect 3775 7040 3781 7104
rect 3845 7040 3861 7104
rect 3925 7040 3941 7104
rect 4005 7040 4021 7104
rect 4085 7040 4091 7104
rect 3775 7039 4091 7040
rect 5661 7104 5977 7105
rect 5661 7040 5667 7104
rect 5731 7040 5747 7104
rect 5811 7040 5827 7104
rect 5891 7040 5907 7104
rect 5971 7040 5977 7104
rect 5661 7039 5977 7040
rect 7547 7104 7863 7105
rect 7547 7040 7553 7104
rect 7617 7040 7633 7104
rect 7697 7040 7713 7104
rect 7777 7040 7793 7104
rect 7857 7040 7863 7104
rect 7547 7039 7863 7040
rect 2549 6560 2865 6561
rect 2549 6496 2555 6560
rect 2619 6496 2635 6560
rect 2699 6496 2715 6560
rect 2779 6496 2795 6560
rect 2859 6496 2865 6560
rect 2549 6495 2865 6496
rect 4435 6560 4751 6561
rect 4435 6496 4441 6560
rect 4505 6496 4521 6560
rect 4585 6496 4601 6560
rect 4665 6496 4681 6560
rect 4745 6496 4751 6560
rect 4435 6495 4751 6496
rect 6321 6560 6637 6561
rect 6321 6496 6327 6560
rect 6391 6496 6407 6560
rect 6471 6496 6487 6560
rect 6551 6496 6567 6560
rect 6631 6496 6637 6560
rect 6321 6495 6637 6496
rect 8207 6560 8523 6561
rect 8207 6496 8213 6560
rect 8277 6496 8293 6560
rect 8357 6496 8373 6560
rect 8437 6496 8453 6560
rect 8517 6496 8523 6560
rect 8207 6495 8523 6496
rect 1889 6016 2205 6017
rect 1889 5952 1895 6016
rect 1959 5952 1975 6016
rect 2039 5952 2055 6016
rect 2119 5952 2135 6016
rect 2199 5952 2205 6016
rect 1889 5951 2205 5952
rect 3775 6016 4091 6017
rect 3775 5952 3781 6016
rect 3845 5952 3861 6016
rect 3925 5952 3941 6016
rect 4005 5952 4021 6016
rect 4085 5952 4091 6016
rect 3775 5951 4091 5952
rect 5661 6016 5977 6017
rect 5661 5952 5667 6016
rect 5731 5952 5747 6016
rect 5811 5952 5827 6016
rect 5891 5952 5907 6016
rect 5971 5952 5977 6016
rect 5661 5951 5977 5952
rect 7547 6016 7863 6017
rect 7547 5952 7553 6016
rect 7617 5952 7633 6016
rect 7697 5952 7713 6016
rect 7777 5952 7793 6016
rect 7857 5952 7863 6016
rect 7547 5951 7863 5952
rect 2549 5472 2865 5473
rect 2549 5408 2555 5472
rect 2619 5408 2635 5472
rect 2699 5408 2715 5472
rect 2779 5408 2795 5472
rect 2859 5408 2865 5472
rect 2549 5407 2865 5408
rect 4435 5472 4751 5473
rect 4435 5408 4441 5472
rect 4505 5408 4521 5472
rect 4585 5408 4601 5472
rect 4665 5408 4681 5472
rect 4745 5408 4751 5472
rect 4435 5407 4751 5408
rect 6321 5472 6637 5473
rect 6321 5408 6327 5472
rect 6391 5408 6407 5472
rect 6471 5408 6487 5472
rect 6551 5408 6567 5472
rect 6631 5408 6637 5472
rect 6321 5407 6637 5408
rect 8207 5472 8523 5473
rect 8207 5408 8213 5472
rect 8277 5408 8293 5472
rect 8357 5408 8373 5472
rect 8437 5408 8453 5472
rect 8517 5408 8523 5472
rect 8207 5407 8523 5408
rect 1889 4928 2205 4929
rect 1889 4864 1895 4928
rect 1959 4864 1975 4928
rect 2039 4864 2055 4928
rect 2119 4864 2135 4928
rect 2199 4864 2205 4928
rect 1889 4863 2205 4864
rect 3775 4928 4091 4929
rect 3775 4864 3781 4928
rect 3845 4864 3861 4928
rect 3925 4864 3941 4928
rect 4005 4864 4021 4928
rect 4085 4864 4091 4928
rect 3775 4863 4091 4864
rect 5661 4928 5977 4929
rect 5661 4864 5667 4928
rect 5731 4864 5747 4928
rect 5811 4864 5827 4928
rect 5891 4864 5907 4928
rect 5971 4864 5977 4928
rect 5661 4863 5977 4864
rect 7547 4928 7863 4929
rect 7547 4864 7553 4928
rect 7617 4864 7633 4928
rect 7697 4864 7713 4928
rect 7777 4864 7793 4928
rect 7857 4864 7863 4928
rect 7547 4863 7863 4864
rect 2549 4384 2865 4385
rect 2549 4320 2555 4384
rect 2619 4320 2635 4384
rect 2699 4320 2715 4384
rect 2779 4320 2795 4384
rect 2859 4320 2865 4384
rect 2549 4319 2865 4320
rect 4435 4384 4751 4385
rect 4435 4320 4441 4384
rect 4505 4320 4521 4384
rect 4585 4320 4601 4384
rect 4665 4320 4681 4384
rect 4745 4320 4751 4384
rect 4435 4319 4751 4320
rect 6321 4384 6637 4385
rect 6321 4320 6327 4384
rect 6391 4320 6407 4384
rect 6471 4320 6487 4384
rect 6551 4320 6567 4384
rect 6631 4320 6637 4384
rect 6321 4319 6637 4320
rect 8207 4384 8523 4385
rect 8207 4320 8213 4384
rect 8277 4320 8293 4384
rect 8357 4320 8373 4384
rect 8437 4320 8453 4384
rect 8517 4320 8523 4384
rect 8207 4319 8523 4320
rect 0 4178 800 4208
rect 1669 4178 1735 4181
rect 0 4176 1735 4178
rect 0 4120 1674 4176
rect 1730 4120 1735 4176
rect 0 4118 1735 4120
rect 0 4088 800 4118
rect 1669 4115 1735 4118
rect 1889 3840 2205 3841
rect 1889 3776 1895 3840
rect 1959 3776 1975 3840
rect 2039 3776 2055 3840
rect 2119 3776 2135 3840
rect 2199 3776 2205 3840
rect 1889 3775 2205 3776
rect 3775 3840 4091 3841
rect 3775 3776 3781 3840
rect 3845 3776 3861 3840
rect 3925 3776 3941 3840
rect 4005 3776 4021 3840
rect 4085 3776 4091 3840
rect 3775 3775 4091 3776
rect 5661 3840 5977 3841
rect 5661 3776 5667 3840
rect 5731 3776 5747 3840
rect 5811 3776 5827 3840
rect 5891 3776 5907 3840
rect 5971 3776 5977 3840
rect 5661 3775 5977 3776
rect 7547 3840 7863 3841
rect 7547 3776 7553 3840
rect 7617 3776 7633 3840
rect 7697 3776 7713 3840
rect 7777 3776 7793 3840
rect 7857 3776 7863 3840
rect 7547 3775 7863 3776
rect 2549 3296 2865 3297
rect 2549 3232 2555 3296
rect 2619 3232 2635 3296
rect 2699 3232 2715 3296
rect 2779 3232 2795 3296
rect 2859 3232 2865 3296
rect 2549 3231 2865 3232
rect 4435 3296 4751 3297
rect 4435 3232 4441 3296
rect 4505 3232 4521 3296
rect 4585 3232 4601 3296
rect 4665 3232 4681 3296
rect 4745 3232 4751 3296
rect 4435 3231 4751 3232
rect 6321 3296 6637 3297
rect 6321 3232 6327 3296
rect 6391 3232 6407 3296
rect 6471 3232 6487 3296
rect 6551 3232 6567 3296
rect 6631 3232 6637 3296
rect 6321 3231 6637 3232
rect 8207 3296 8523 3297
rect 8207 3232 8213 3296
rect 8277 3232 8293 3296
rect 8357 3232 8373 3296
rect 8437 3232 8453 3296
rect 8517 3232 8523 3296
rect 8207 3231 8523 3232
rect 8017 2818 8083 2821
rect 8978 2818 9778 2848
rect 8017 2816 9778 2818
rect 8017 2760 8022 2816
rect 8078 2760 9778 2816
rect 8017 2758 9778 2760
rect 8017 2755 8083 2758
rect 1889 2752 2205 2753
rect 1889 2688 1895 2752
rect 1959 2688 1975 2752
rect 2039 2688 2055 2752
rect 2119 2688 2135 2752
rect 2199 2688 2205 2752
rect 1889 2687 2205 2688
rect 3775 2752 4091 2753
rect 3775 2688 3781 2752
rect 3845 2688 3861 2752
rect 3925 2688 3941 2752
rect 4005 2688 4021 2752
rect 4085 2688 4091 2752
rect 3775 2687 4091 2688
rect 5661 2752 5977 2753
rect 5661 2688 5667 2752
rect 5731 2688 5747 2752
rect 5811 2688 5827 2752
rect 5891 2688 5907 2752
rect 5971 2688 5977 2752
rect 5661 2687 5977 2688
rect 7547 2752 7863 2753
rect 7547 2688 7553 2752
rect 7617 2688 7633 2752
rect 7697 2688 7713 2752
rect 7777 2688 7793 2752
rect 7857 2688 7863 2752
rect 8978 2728 9778 2758
rect 7547 2687 7863 2688
rect 2549 2208 2865 2209
rect 2549 2144 2555 2208
rect 2619 2144 2635 2208
rect 2699 2144 2715 2208
rect 2779 2144 2795 2208
rect 2859 2144 2865 2208
rect 2549 2143 2865 2144
rect 4435 2208 4751 2209
rect 4435 2144 4441 2208
rect 4505 2144 4521 2208
rect 4585 2144 4601 2208
rect 4665 2144 4681 2208
rect 4745 2144 4751 2208
rect 4435 2143 4751 2144
rect 6321 2208 6637 2209
rect 6321 2144 6327 2208
rect 6391 2144 6407 2208
rect 6471 2144 6487 2208
rect 6551 2144 6567 2208
rect 6631 2144 6637 2208
rect 6321 2143 6637 2144
rect 8207 2208 8523 2209
rect 8207 2144 8213 2208
rect 8277 2144 8293 2208
rect 8357 2144 8373 2208
rect 8437 2144 8453 2208
rect 8517 2144 8523 2208
rect 8207 2143 8523 2144
<< via3 >>
rect 1895 9276 1959 9280
rect 1895 9220 1899 9276
rect 1899 9220 1955 9276
rect 1955 9220 1959 9276
rect 1895 9216 1959 9220
rect 1975 9276 2039 9280
rect 1975 9220 1979 9276
rect 1979 9220 2035 9276
rect 2035 9220 2039 9276
rect 1975 9216 2039 9220
rect 2055 9276 2119 9280
rect 2055 9220 2059 9276
rect 2059 9220 2115 9276
rect 2115 9220 2119 9276
rect 2055 9216 2119 9220
rect 2135 9276 2199 9280
rect 2135 9220 2139 9276
rect 2139 9220 2195 9276
rect 2195 9220 2199 9276
rect 2135 9216 2199 9220
rect 3781 9276 3845 9280
rect 3781 9220 3785 9276
rect 3785 9220 3841 9276
rect 3841 9220 3845 9276
rect 3781 9216 3845 9220
rect 3861 9276 3925 9280
rect 3861 9220 3865 9276
rect 3865 9220 3921 9276
rect 3921 9220 3925 9276
rect 3861 9216 3925 9220
rect 3941 9276 4005 9280
rect 3941 9220 3945 9276
rect 3945 9220 4001 9276
rect 4001 9220 4005 9276
rect 3941 9216 4005 9220
rect 4021 9276 4085 9280
rect 4021 9220 4025 9276
rect 4025 9220 4081 9276
rect 4081 9220 4085 9276
rect 4021 9216 4085 9220
rect 5667 9276 5731 9280
rect 5667 9220 5671 9276
rect 5671 9220 5727 9276
rect 5727 9220 5731 9276
rect 5667 9216 5731 9220
rect 5747 9276 5811 9280
rect 5747 9220 5751 9276
rect 5751 9220 5807 9276
rect 5807 9220 5811 9276
rect 5747 9216 5811 9220
rect 5827 9276 5891 9280
rect 5827 9220 5831 9276
rect 5831 9220 5887 9276
rect 5887 9220 5891 9276
rect 5827 9216 5891 9220
rect 5907 9276 5971 9280
rect 5907 9220 5911 9276
rect 5911 9220 5967 9276
rect 5967 9220 5971 9276
rect 5907 9216 5971 9220
rect 7553 9276 7617 9280
rect 7553 9220 7557 9276
rect 7557 9220 7613 9276
rect 7613 9220 7617 9276
rect 7553 9216 7617 9220
rect 7633 9276 7697 9280
rect 7633 9220 7637 9276
rect 7637 9220 7693 9276
rect 7693 9220 7697 9276
rect 7633 9216 7697 9220
rect 7713 9276 7777 9280
rect 7713 9220 7717 9276
rect 7717 9220 7773 9276
rect 7773 9220 7777 9276
rect 7713 9216 7777 9220
rect 7793 9276 7857 9280
rect 7793 9220 7797 9276
rect 7797 9220 7853 9276
rect 7853 9220 7857 9276
rect 7793 9216 7857 9220
rect 2555 8732 2619 8736
rect 2555 8676 2559 8732
rect 2559 8676 2615 8732
rect 2615 8676 2619 8732
rect 2555 8672 2619 8676
rect 2635 8732 2699 8736
rect 2635 8676 2639 8732
rect 2639 8676 2695 8732
rect 2695 8676 2699 8732
rect 2635 8672 2699 8676
rect 2715 8732 2779 8736
rect 2715 8676 2719 8732
rect 2719 8676 2775 8732
rect 2775 8676 2779 8732
rect 2715 8672 2779 8676
rect 2795 8732 2859 8736
rect 2795 8676 2799 8732
rect 2799 8676 2855 8732
rect 2855 8676 2859 8732
rect 2795 8672 2859 8676
rect 4441 8732 4505 8736
rect 4441 8676 4445 8732
rect 4445 8676 4501 8732
rect 4501 8676 4505 8732
rect 4441 8672 4505 8676
rect 4521 8732 4585 8736
rect 4521 8676 4525 8732
rect 4525 8676 4581 8732
rect 4581 8676 4585 8732
rect 4521 8672 4585 8676
rect 4601 8732 4665 8736
rect 4601 8676 4605 8732
rect 4605 8676 4661 8732
rect 4661 8676 4665 8732
rect 4601 8672 4665 8676
rect 4681 8732 4745 8736
rect 4681 8676 4685 8732
rect 4685 8676 4741 8732
rect 4741 8676 4745 8732
rect 4681 8672 4745 8676
rect 6327 8732 6391 8736
rect 6327 8676 6331 8732
rect 6331 8676 6387 8732
rect 6387 8676 6391 8732
rect 6327 8672 6391 8676
rect 6407 8732 6471 8736
rect 6407 8676 6411 8732
rect 6411 8676 6467 8732
rect 6467 8676 6471 8732
rect 6407 8672 6471 8676
rect 6487 8732 6551 8736
rect 6487 8676 6491 8732
rect 6491 8676 6547 8732
rect 6547 8676 6551 8732
rect 6487 8672 6551 8676
rect 6567 8732 6631 8736
rect 6567 8676 6571 8732
rect 6571 8676 6627 8732
rect 6627 8676 6631 8732
rect 6567 8672 6631 8676
rect 8213 8732 8277 8736
rect 8213 8676 8217 8732
rect 8217 8676 8273 8732
rect 8273 8676 8277 8732
rect 8213 8672 8277 8676
rect 8293 8732 8357 8736
rect 8293 8676 8297 8732
rect 8297 8676 8353 8732
rect 8353 8676 8357 8732
rect 8293 8672 8357 8676
rect 8373 8732 8437 8736
rect 8373 8676 8377 8732
rect 8377 8676 8433 8732
rect 8433 8676 8437 8732
rect 8373 8672 8437 8676
rect 8453 8732 8517 8736
rect 8453 8676 8457 8732
rect 8457 8676 8513 8732
rect 8513 8676 8517 8732
rect 8453 8672 8517 8676
rect 1895 8188 1959 8192
rect 1895 8132 1899 8188
rect 1899 8132 1955 8188
rect 1955 8132 1959 8188
rect 1895 8128 1959 8132
rect 1975 8188 2039 8192
rect 1975 8132 1979 8188
rect 1979 8132 2035 8188
rect 2035 8132 2039 8188
rect 1975 8128 2039 8132
rect 2055 8188 2119 8192
rect 2055 8132 2059 8188
rect 2059 8132 2115 8188
rect 2115 8132 2119 8188
rect 2055 8128 2119 8132
rect 2135 8188 2199 8192
rect 2135 8132 2139 8188
rect 2139 8132 2195 8188
rect 2195 8132 2199 8188
rect 2135 8128 2199 8132
rect 3781 8188 3845 8192
rect 3781 8132 3785 8188
rect 3785 8132 3841 8188
rect 3841 8132 3845 8188
rect 3781 8128 3845 8132
rect 3861 8188 3925 8192
rect 3861 8132 3865 8188
rect 3865 8132 3921 8188
rect 3921 8132 3925 8188
rect 3861 8128 3925 8132
rect 3941 8188 4005 8192
rect 3941 8132 3945 8188
rect 3945 8132 4001 8188
rect 4001 8132 4005 8188
rect 3941 8128 4005 8132
rect 4021 8188 4085 8192
rect 4021 8132 4025 8188
rect 4025 8132 4081 8188
rect 4081 8132 4085 8188
rect 4021 8128 4085 8132
rect 5667 8188 5731 8192
rect 5667 8132 5671 8188
rect 5671 8132 5727 8188
rect 5727 8132 5731 8188
rect 5667 8128 5731 8132
rect 5747 8188 5811 8192
rect 5747 8132 5751 8188
rect 5751 8132 5807 8188
rect 5807 8132 5811 8188
rect 5747 8128 5811 8132
rect 5827 8188 5891 8192
rect 5827 8132 5831 8188
rect 5831 8132 5887 8188
rect 5887 8132 5891 8188
rect 5827 8128 5891 8132
rect 5907 8188 5971 8192
rect 5907 8132 5911 8188
rect 5911 8132 5967 8188
rect 5967 8132 5971 8188
rect 5907 8128 5971 8132
rect 7553 8188 7617 8192
rect 7553 8132 7557 8188
rect 7557 8132 7613 8188
rect 7613 8132 7617 8188
rect 7553 8128 7617 8132
rect 7633 8188 7697 8192
rect 7633 8132 7637 8188
rect 7637 8132 7693 8188
rect 7693 8132 7697 8188
rect 7633 8128 7697 8132
rect 7713 8188 7777 8192
rect 7713 8132 7717 8188
rect 7717 8132 7773 8188
rect 7773 8132 7777 8188
rect 7713 8128 7777 8132
rect 7793 8188 7857 8192
rect 7793 8132 7797 8188
rect 7797 8132 7853 8188
rect 7853 8132 7857 8188
rect 7793 8128 7857 8132
rect 2555 7644 2619 7648
rect 2555 7588 2559 7644
rect 2559 7588 2615 7644
rect 2615 7588 2619 7644
rect 2555 7584 2619 7588
rect 2635 7644 2699 7648
rect 2635 7588 2639 7644
rect 2639 7588 2695 7644
rect 2695 7588 2699 7644
rect 2635 7584 2699 7588
rect 2715 7644 2779 7648
rect 2715 7588 2719 7644
rect 2719 7588 2775 7644
rect 2775 7588 2779 7644
rect 2715 7584 2779 7588
rect 2795 7644 2859 7648
rect 2795 7588 2799 7644
rect 2799 7588 2855 7644
rect 2855 7588 2859 7644
rect 2795 7584 2859 7588
rect 4441 7644 4505 7648
rect 4441 7588 4445 7644
rect 4445 7588 4501 7644
rect 4501 7588 4505 7644
rect 4441 7584 4505 7588
rect 4521 7644 4585 7648
rect 4521 7588 4525 7644
rect 4525 7588 4581 7644
rect 4581 7588 4585 7644
rect 4521 7584 4585 7588
rect 4601 7644 4665 7648
rect 4601 7588 4605 7644
rect 4605 7588 4661 7644
rect 4661 7588 4665 7644
rect 4601 7584 4665 7588
rect 4681 7644 4745 7648
rect 4681 7588 4685 7644
rect 4685 7588 4741 7644
rect 4741 7588 4745 7644
rect 4681 7584 4745 7588
rect 6327 7644 6391 7648
rect 6327 7588 6331 7644
rect 6331 7588 6387 7644
rect 6387 7588 6391 7644
rect 6327 7584 6391 7588
rect 6407 7644 6471 7648
rect 6407 7588 6411 7644
rect 6411 7588 6467 7644
rect 6467 7588 6471 7644
rect 6407 7584 6471 7588
rect 6487 7644 6551 7648
rect 6487 7588 6491 7644
rect 6491 7588 6547 7644
rect 6547 7588 6551 7644
rect 6487 7584 6551 7588
rect 6567 7644 6631 7648
rect 6567 7588 6571 7644
rect 6571 7588 6627 7644
rect 6627 7588 6631 7644
rect 6567 7584 6631 7588
rect 8213 7644 8277 7648
rect 8213 7588 8217 7644
rect 8217 7588 8273 7644
rect 8273 7588 8277 7644
rect 8213 7584 8277 7588
rect 8293 7644 8357 7648
rect 8293 7588 8297 7644
rect 8297 7588 8353 7644
rect 8353 7588 8357 7644
rect 8293 7584 8357 7588
rect 8373 7644 8437 7648
rect 8373 7588 8377 7644
rect 8377 7588 8433 7644
rect 8433 7588 8437 7644
rect 8373 7584 8437 7588
rect 8453 7644 8517 7648
rect 8453 7588 8457 7644
rect 8457 7588 8513 7644
rect 8513 7588 8517 7644
rect 8453 7584 8517 7588
rect 1895 7100 1959 7104
rect 1895 7044 1899 7100
rect 1899 7044 1955 7100
rect 1955 7044 1959 7100
rect 1895 7040 1959 7044
rect 1975 7100 2039 7104
rect 1975 7044 1979 7100
rect 1979 7044 2035 7100
rect 2035 7044 2039 7100
rect 1975 7040 2039 7044
rect 2055 7100 2119 7104
rect 2055 7044 2059 7100
rect 2059 7044 2115 7100
rect 2115 7044 2119 7100
rect 2055 7040 2119 7044
rect 2135 7100 2199 7104
rect 2135 7044 2139 7100
rect 2139 7044 2195 7100
rect 2195 7044 2199 7100
rect 2135 7040 2199 7044
rect 3781 7100 3845 7104
rect 3781 7044 3785 7100
rect 3785 7044 3841 7100
rect 3841 7044 3845 7100
rect 3781 7040 3845 7044
rect 3861 7100 3925 7104
rect 3861 7044 3865 7100
rect 3865 7044 3921 7100
rect 3921 7044 3925 7100
rect 3861 7040 3925 7044
rect 3941 7100 4005 7104
rect 3941 7044 3945 7100
rect 3945 7044 4001 7100
rect 4001 7044 4005 7100
rect 3941 7040 4005 7044
rect 4021 7100 4085 7104
rect 4021 7044 4025 7100
rect 4025 7044 4081 7100
rect 4081 7044 4085 7100
rect 4021 7040 4085 7044
rect 5667 7100 5731 7104
rect 5667 7044 5671 7100
rect 5671 7044 5727 7100
rect 5727 7044 5731 7100
rect 5667 7040 5731 7044
rect 5747 7100 5811 7104
rect 5747 7044 5751 7100
rect 5751 7044 5807 7100
rect 5807 7044 5811 7100
rect 5747 7040 5811 7044
rect 5827 7100 5891 7104
rect 5827 7044 5831 7100
rect 5831 7044 5887 7100
rect 5887 7044 5891 7100
rect 5827 7040 5891 7044
rect 5907 7100 5971 7104
rect 5907 7044 5911 7100
rect 5911 7044 5967 7100
rect 5967 7044 5971 7100
rect 5907 7040 5971 7044
rect 7553 7100 7617 7104
rect 7553 7044 7557 7100
rect 7557 7044 7613 7100
rect 7613 7044 7617 7100
rect 7553 7040 7617 7044
rect 7633 7100 7697 7104
rect 7633 7044 7637 7100
rect 7637 7044 7693 7100
rect 7693 7044 7697 7100
rect 7633 7040 7697 7044
rect 7713 7100 7777 7104
rect 7713 7044 7717 7100
rect 7717 7044 7773 7100
rect 7773 7044 7777 7100
rect 7713 7040 7777 7044
rect 7793 7100 7857 7104
rect 7793 7044 7797 7100
rect 7797 7044 7853 7100
rect 7853 7044 7857 7100
rect 7793 7040 7857 7044
rect 2555 6556 2619 6560
rect 2555 6500 2559 6556
rect 2559 6500 2615 6556
rect 2615 6500 2619 6556
rect 2555 6496 2619 6500
rect 2635 6556 2699 6560
rect 2635 6500 2639 6556
rect 2639 6500 2695 6556
rect 2695 6500 2699 6556
rect 2635 6496 2699 6500
rect 2715 6556 2779 6560
rect 2715 6500 2719 6556
rect 2719 6500 2775 6556
rect 2775 6500 2779 6556
rect 2715 6496 2779 6500
rect 2795 6556 2859 6560
rect 2795 6500 2799 6556
rect 2799 6500 2855 6556
rect 2855 6500 2859 6556
rect 2795 6496 2859 6500
rect 4441 6556 4505 6560
rect 4441 6500 4445 6556
rect 4445 6500 4501 6556
rect 4501 6500 4505 6556
rect 4441 6496 4505 6500
rect 4521 6556 4585 6560
rect 4521 6500 4525 6556
rect 4525 6500 4581 6556
rect 4581 6500 4585 6556
rect 4521 6496 4585 6500
rect 4601 6556 4665 6560
rect 4601 6500 4605 6556
rect 4605 6500 4661 6556
rect 4661 6500 4665 6556
rect 4601 6496 4665 6500
rect 4681 6556 4745 6560
rect 4681 6500 4685 6556
rect 4685 6500 4741 6556
rect 4741 6500 4745 6556
rect 4681 6496 4745 6500
rect 6327 6556 6391 6560
rect 6327 6500 6331 6556
rect 6331 6500 6387 6556
rect 6387 6500 6391 6556
rect 6327 6496 6391 6500
rect 6407 6556 6471 6560
rect 6407 6500 6411 6556
rect 6411 6500 6467 6556
rect 6467 6500 6471 6556
rect 6407 6496 6471 6500
rect 6487 6556 6551 6560
rect 6487 6500 6491 6556
rect 6491 6500 6547 6556
rect 6547 6500 6551 6556
rect 6487 6496 6551 6500
rect 6567 6556 6631 6560
rect 6567 6500 6571 6556
rect 6571 6500 6627 6556
rect 6627 6500 6631 6556
rect 6567 6496 6631 6500
rect 8213 6556 8277 6560
rect 8213 6500 8217 6556
rect 8217 6500 8273 6556
rect 8273 6500 8277 6556
rect 8213 6496 8277 6500
rect 8293 6556 8357 6560
rect 8293 6500 8297 6556
rect 8297 6500 8353 6556
rect 8353 6500 8357 6556
rect 8293 6496 8357 6500
rect 8373 6556 8437 6560
rect 8373 6500 8377 6556
rect 8377 6500 8433 6556
rect 8433 6500 8437 6556
rect 8373 6496 8437 6500
rect 8453 6556 8517 6560
rect 8453 6500 8457 6556
rect 8457 6500 8513 6556
rect 8513 6500 8517 6556
rect 8453 6496 8517 6500
rect 1895 6012 1959 6016
rect 1895 5956 1899 6012
rect 1899 5956 1955 6012
rect 1955 5956 1959 6012
rect 1895 5952 1959 5956
rect 1975 6012 2039 6016
rect 1975 5956 1979 6012
rect 1979 5956 2035 6012
rect 2035 5956 2039 6012
rect 1975 5952 2039 5956
rect 2055 6012 2119 6016
rect 2055 5956 2059 6012
rect 2059 5956 2115 6012
rect 2115 5956 2119 6012
rect 2055 5952 2119 5956
rect 2135 6012 2199 6016
rect 2135 5956 2139 6012
rect 2139 5956 2195 6012
rect 2195 5956 2199 6012
rect 2135 5952 2199 5956
rect 3781 6012 3845 6016
rect 3781 5956 3785 6012
rect 3785 5956 3841 6012
rect 3841 5956 3845 6012
rect 3781 5952 3845 5956
rect 3861 6012 3925 6016
rect 3861 5956 3865 6012
rect 3865 5956 3921 6012
rect 3921 5956 3925 6012
rect 3861 5952 3925 5956
rect 3941 6012 4005 6016
rect 3941 5956 3945 6012
rect 3945 5956 4001 6012
rect 4001 5956 4005 6012
rect 3941 5952 4005 5956
rect 4021 6012 4085 6016
rect 4021 5956 4025 6012
rect 4025 5956 4081 6012
rect 4081 5956 4085 6012
rect 4021 5952 4085 5956
rect 5667 6012 5731 6016
rect 5667 5956 5671 6012
rect 5671 5956 5727 6012
rect 5727 5956 5731 6012
rect 5667 5952 5731 5956
rect 5747 6012 5811 6016
rect 5747 5956 5751 6012
rect 5751 5956 5807 6012
rect 5807 5956 5811 6012
rect 5747 5952 5811 5956
rect 5827 6012 5891 6016
rect 5827 5956 5831 6012
rect 5831 5956 5887 6012
rect 5887 5956 5891 6012
rect 5827 5952 5891 5956
rect 5907 6012 5971 6016
rect 5907 5956 5911 6012
rect 5911 5956 5967 6012
rect 5967 5956 5971 6012
rect 5907 5952 5971 5956
rect 7553 6012 7617 6016
rect 7553 5956 7557 6012
rect 7557 5956 7613 6012
rect 7613 5956 7617 6012
rect 7553 5952 7617 5956
rect 7633 6012 7697 6016
rect 7633 5956 7637 6012
rect 7637 5956 7693 6012
rect 7693 5956 7697 6012
rect 7633 5952 7697 5956
rect 7713 6012 7777 6016
rect 7713 5956 7717 6012
rect 7717 5956 7773 6012
rect 7773 5956 7777 6012
rect 7713 5952 7777 5956
rect 7793 6012 7857 6016
rect 7793 5956 7797 6012
rect 7797 5956 7853 6012
rect 7853 5956 7857 6012
rect 7793 5952 7857 5956
rect 2555 5468 2619 5472
rect 2555 5412 2559 5468
rect 2559 5412 2615 5468
rect 2615 5412 2619 5468
rect 2555 5408 2619 5412
rect 2635 5468 2699 5472
rect 2635 5412 2639 5468
rect 2639 5412 2695 5468
rect 2695 5412 2699 5468
rect 2635 5408 2699 5412
rect 2715 5468 2779 5472
rect 2715 5412 2719 5468
rect 2719 5412 2775 5468
rect 2775 5412 2779 5468
rect 2715 5408 2779 5412
rect 2795 5468 2859 5472
rect 2795 5412 2799 5468
rect 2799 5412 2855 5468
rect 2855 5412 2859 5468
rect 2795 5408 2859 5412
rect 4441 5468 4505 5472
rect 4441 5412 4445 5468
rect 4445 5412 4501 5468
rect 4501 5412 4505 5468
rect 4441 5408 4505 5412
rect 4521 5468 4585 5472
rect 4521 5412 4525 5468
rect 4525 5412 4581 5468
rect 4581 5412 4585 5468
rect 4521 5408 4585 5412
rect 4601 5468 4665 5472
rect 4601 5412 4605 5468
rect 4605 5412 4661 5468
rect 4661 5412 4665 5468
rect 4601 5408 4665 5412
rect 4681 5468 4745 5472
rect 4681 5412 4685 5468
rect 4685 5412 4741 5468
rect 4741 5412 4745 5468
rect 4681 5408 4745 5412
rect 6327 5468 6391 5472
rect 6327 5412 6331 5468
rect 6331 5412 6387 5468
rect 6387 5412 6391 5468
rect 6327 5408 6391 5412
rect 6407 5468 6471 5472
rect 6407 5412 6411 5468
rect 6411 5412 6467 5468
rect 6467 5412 6471 5468
rect 6407 5408 6471 5412
rect 6487 5468 6551 5472
rect 6487 5412 6491 5468
rect 6491 5412 6547 5468
rect 6547 5412 6551 5468
rect 6487 5408 6551 5412
rect 6567 5468 6631 5472
rect 6567 5412 6571 5468
rect 6571 5412 6627 5468
rect 6627 5412 6631 5468
rect 6567 5408 6631 5412
rect 8213 5468 8277 5472
rect 8213 5412 8217 5468
rect 8217 5412 8273 5468
rect 8273 5412 8277 5468
rect 8213 5408 8277 5412
rect 8293 5468 8357 5472
rect 8293 5412 8297 5468
rect 8297 5412 8353 5468
rect 8353 5412 8357 5468
rect 8293 5408 8357 5412
rect 8373 5468 8437 5472
rect 8373 5412 8377 5468
rect 8377 5412 8433 5468
rect 8433 5412 8437 5468
rect 8373 5408 8437 5412
rect 8453 5468 8517 5472
rect 8453 5412 8457 5468
rect 8457 5412 8513 5468
rect 8513 5412 8517 5468
rect 8453 5408 8517 5412
rect 1895 4924 1959 4928
rect 1895 4868 1899 4924
rect 1899 4868 1955 4924
rect 1955 4868 1959 4924
rect 1895 4864 1959 4868
rect 1975 4924 2039 4928
rect 1975 4868 1979 4924
rect 1979 4868 2035 4924
rect 2035 4868 2039 4924
rect 1975 4864 2039 4868
rect 2055 4924 2119 4928
rect 2055 4868 2059 4924
rect 2059 4868 2115 4924
rect 2115 4868 2119 4924
rect 2055 4864 2119 4868
rect 2135 4924 2199 4928
rect 2135 4868 2139 4924
rect 2139 4868 2195 4924
rect 2195 4868 2199 4924
rect 2135 4864 2199 4868
rect 3781 4924 3845 4928
rect 3781 4868 3785 4924
rect 3785 4868 3841 4924
rect 3841 4868 3845 4924
rect 3781 4864 3845 4868
rect 3861 4924 3925 4928
rect 3861 4868 3865 4924
rect 3865 4868 3921 4924
rect 3921 4868 3925 4924
rect 3861 4864 3925 4868
rect 3941 4924 4005 4928
rect 3941 4868 3945 4924
rect 3945 4868 4001 4924
rect 4001 4868 4005 4924
rect 3941 4864 4005 4868
rect 4021 4924 4085 4928
rect 4021 4868 4025 4924
rect 4025 4868 4081 4924
rect 4081 4868 4085 4924
rect 4021 4864 4085 4868
rect 5667 4924 5731 4928
rect 5667 4868 5671 4924
rect 5671 4868 5727 4924
rect 5727 4868 5731 4924
rect 5667 4864 5731 4868
rect 5747 4924 5811 4928
rect 5747 4868 5751 4924
rect 5751 4868 5807 4924
rect 5807 4868 5811 4924
rect 5747 4864 5811 4868
rect 5827 4924 5891 4928
rect 5827 4868 5831 4924
rect 5831 4868 5887 4924
rect 5887 4868 5891 4924
rect 5827 4864 5891 4868
rect 5907 4924 5971 4928
rect 5907 4868 5911 4924
rect 5911 4868 5967 4924
rect 5967 4868 5971 4924
rect 5907 4864 5971 4868
rect 7553 4924 7617 4928
rect 7553 4868 7557 4924
rect 7557 4868 7613 4924
rect 7613 4868 7617 4924
rect 7553 4864 7617 4868
rect 7633 4924 7697 4928
rect 7633 4868 7637 4924
rect 7637 4868 7693 4924
rect 7693 4868 7697 4924
rect 7633 4864 7697 4868
rect 7713 4924 7777 4928
rect 7713 4868 7717 4924
rect 7717 4868 7773 4924
rect 7773 4868 7777 4924
rect 7713 4864 7777 4868
rect 7793 4924 7857 4928
rect 7793 4868 7797 4924
rect 7797 4868 7853 4924
rect 7853 4868 7857 4924
rect 7793 4864 7857 4868
rect 2555 4380 2619 4384
rect 2555 4324 2559 4380
rect 2559 4324 2615 4380
rect 2615 4324 2619 4380
rect 2555 4320 2619 4324
rect 2635 4380 2699 4384
rect 2635 4324 2639 4380
rect 2639 4324 2695 4380
rect 2695 4324 2699 4380
rect 2635 4320 2699 4324
rect 2715 4380 2779 4384
rect 2715 4324 2719 4380
rect 2719 4324 2775 4380
rect 2775 4324 2779 4380
rect 2715 4320 2779 4324
rect 2795 4380 2859 4384
rect 2795 4324 2799 4380
rect 2799 4324 2855 4380
rect 2855 4324 2859 4380
rect 2795 4320 2859 4324
rect 4441 4380 4505 4384
rect 4441 4324 4445 4380
rect 4445 4324 4501 4380
rect 4501 4324 4505 4380
rect 4441 4320 4505 4324
rect 4521 4380 4585 4384
rect 4521 4324 4525 4380
rect 4525 4324 4581 4380
rect 4581 4324 4585 4380
rect 4521 4320 4585 4324
rect 4601 4380 4665 4384
rect 4601 4324 4605 4380
rect 4605 4324 4661 4380
rect 4661 4324 4665 4380
rect 4601 4320 4665 4324
rect 4681 4380 4745 4384
rect 4681 4324 4685 4380
rect 4685 4324 4741 4380
rect 4741 4324 4745 4380
rect 4681 4320 4745 4324
rect 6327 4380 6391 4384
rect 6327 4324 6331 4380
rect 6331 4324 6387 4380
rect 6387 4324 6391 4380
rect 6327 4320 6391 4324
rect 6407 4380 6471 4384
rect 6407 4324 6411 4380
rect 6411 4324 6467 4380
rect 6467 4324 6471 4380
rect 6407 4320 6471 4324
rect 6487 4380 6551 4384
rect 6487 4324 6491 4380
rect 6491 4324 6547 4380
rect 6547 4324 6551 4380
rect 6487 4320 6551 4324
rect 6567 4380 6631 4384
rect 6567 4324 6571 4380
rect 6571 4324 6627 4380
rect 6627 4324 6631 4380
rect 6567 4320 6631 4324
rect 8213 4380 8277 4384
rect 8213 4324 8217 4380
rect 8217 4324 8273 4380
rect 8273 4324 8277 4380
rect 8213 4320 8277 4324
rect 8293 4380 8357 4384
rect 8293 4324 8297 4380
rect 8297 4324 8353 4380
rect 8353 4324 8357 4380
rect 8293 4320 8357 4324
rect 8373 4380 8437 4384
rect 8373 4324 8377 4380
rect 8377 4324 8433 4380
rect 8433 4324 8437 4380
rect 8373 4320 8437 4324
rect 8453 4380 8517 4384
rect 8453 4324 8457 4380
rect 8457 4324 8513 4380
rect 8513 4324 8517 4380
rect 8453 4320 8517 4324
rect 1895 3836 1959 3840
rect 1895 3780 1899 3836
rect 1899 3780 1955 3836
rect 1955 3780 1959 3836
rect 1895 3776 1959 3780
rect 1975 3836 2039 3840
rect 1975 3780 1979 3836
rect 1979 3780 2035 3836
rect 2035 3780 2039 3836
rect 1975 3776 2039 3780
rect 2055 3836 2119 3840
rect 2055 3780 2059 3836
rect 2059 3780 2115 3836
rect 2115 3780 2119 3836
rect 2055 3776 2119 3780
rect 2135 3836 2199 3840
rect 2135 3780 2139 3836
rect 2139 3780 2195 3836
rect 2195 3780 2199 3836
rect 2135 3776 2199 3780
rect 3781 3836 3845 3840
rect 3781 3780 3785 3836
rect 3785 3780 3841 3836
rect 3841 3780 3845 3836
rect 3781 3776 3845 3780
rect 3861 3836 3925 3840
rect 3861 3780 3865 3836
rect 3865 3780 3921 3836
rect 3921 3780 3925 3836
rect 3861 3776 3925 3780
rect 3941 3836 4005 3840
rect 3941 3780 3945 3836
rect 3945 3780 4001 3836
rect 4001 3780 4005 3836
rect 3941 3776 4005 3780
rect 4021 3836 4085 3840
rect 4021 3780 4025 3836
rect 4025 3780 4081 3836
rect 4081 3780 4085 3836
rect 4021 3776 4085 3780
rect 5667 3836 5731 3840
rect 5667 3780 5671 3836
rect 5671 3780 5727 3836
rect 5727 3780 5731 3836
rect 5667 3776 5731 3780
rect 5747 3836 5811 3840
rect 5747 3780 5751 3836
rect 5751 3780 5807 3836
rect 5807 3780 5811 3836
rect 5747 3776 5811 3780
rect 5827 3836 5891 3840
rect 5827 3780 5831 3836
rect 5831 3780 5887 3836
rect 5887 3780 5891 3836
rect 5827 3776 5891 3780
rect 5907 3836 5971 3840
rect 5907 3780 5911 3836
rect 5911 3780 5967 3836
rect 5967 3780 5971 3836
rect 5907 3776 5971 3780
rect 7553 3836 7617 3840
rect 7553 3780 7557 3836
rect 7557 3780 7613 3836
rect 7613 3780 7617 3836
rect 7553 3776 7617 3780
rect 7633 3836 7697 3840
rect 7633 3780 7637 3836
rect 7637 3780 7693 3836
rect 7693 3780 7697 3836
rect 7633 3776 7697 3780
rect 7713 3836 7777 3840
rect 7713 3780 7717 3836
rect 7717 3780 7773 3836
rect 7773 3780 7777 3836
rect 7713 3776 7777 3780
rect 7793 3836 7857 3840
rect 7793 3780 7797 3836
rect 7797 3780 7853 3836
rect 7853 3780 7857 3836
rect 7793 3776 7857 3780
rect 2555 3292 2619 3296
rect 2555 3236 2559 3292
rect 2559 3236 2615 3292
rect 2615 3236 2619 3292
rect 2555 3232 2619 3236
rect 2635 3292 2699 3296
rect 2635 3236 2639 3292
rect 2639 3236 2695 3292
rect 2695 3236 2699 3292
rect 2635 3232 2699 3236
rect 2715 3292 2779 3296
rect 2715 3236 2719 3292
rect 2719 3236 2775 3292
rect 2775 3236 2779 3292
rect 2715 3232 2779 3236
rect 2795 3292 2859 3296
rect 2795 3236 2799 3292
rect 2799 3236 2855 3292
rect 2855 3236 2859 3292
rect 2795 3232 2859 3236
rect 4441 3292 4505 3296
rect 4441 3236 4445 3292
rect 4445 3236 4501 3292
rect 4501 3236 4505 3292
rect 4441 3232 4505 3236
rect 4521 3292 4585 3296
rect 4521 3236 4525 3292
rect 4525 3236 4581 3292
rect 4581 3236 4585 3292
rect 4521 3232 4585 3236
rect 4601 3292 4665 3296
rect 4601 3236 4605 3292
rect 4605 3236 4661 3292
rect 4661 3236 4665 3292
rect 4601 3232 4665 3236
rect 4681 3292 4745 3296
rect 4681 3236 4685 3292
rect 4685 3236 4741 3292
rect 4741 3236 4745 3292
rect 4681 3232 4745 3236
rect 6327 3292 6391 3296
rect 6327 3236 6331 3292
rect 6331 3236 6387 3292
rect 6387 3236 6391 3292
rect 6327 3232 6391 3236
rect 6407 3292 6471 3296
rect 6407 3236 6411 3292
rect 6411 3236 6467 3292
rect 6467 3236 6471 3292
rect 6407 3232 6471 3236
rect 6487 3292 6551 3296
rect 6487 3236 6491 3292
rect 6491 3236 6547 3292
rect 6547 3236 6551 3292
rect 6487 3232 6551 3236
rect 6567 3292 6631 3296
rect 6567 3236 6571 3292
rect 6571 3236 6627 3292
rect 6627 3236 6631 3292
rect 6567 3232 6631 3236
rect 8213 3292 8277 3296
rect 8213 3236 8217 3292
rect 8217 3236 8273 3292
rect 8273 3236 8277 3292
rect 8213 3232 8277 3236
rect 8293 3292 8357 3296
rect 8293 3236 8297 3292
rect 8297 3236 8353 3292
rect 8353 3236 8357 3292
rect 8293 3232 8357 3236
rect 8373 3292 8437 3296
rect 8373 3236 8377 3292
rect 8377 3236 8433 3292
rect 8433 3236 8437 3292
rect 8373 3232 8437 3236
rect 8453 3292 8517 3296
rect 8453 3236 8457 3292
rect 8457 3236 8513 3292
rect 8513 3236 8517 3292
rect 8453 3232 8517 3236
rect 1895 2748 1959 2752
rect 1895 2692 1899 2748
rect 1899 2692 1955 2748
rect 1955 2692 1959 2748
rect 1895 2688 1959 2692
rect 1975 2748 2039 2752
rect 1975 2692 1979 2748
rect 1979 2692 2035 2748
rect 2035 2692 2039 2748
rect 1975 2688 2039 2692
rect 2055 2748 2119 2752
rect 2055 2692 2059 2748
rect 2059 2692 2115 2748
rect 2115 2692 2119 2748
rect 2055 2688 2119 2692
rect 2135 2748 2199 2752
rect 2135 2692 2139 2748
rect 2139 2692 2195 2748
rect 2195 2692 2199 2748
rect 2135 2688 2199 2692
rect 3781 2748 3845 2752
rect 3781 2692 3785 2748
rect 3785 2692 3841 2748
rect 3841 2692 3845 2748
rect 3781 2688 3845 2692
rect 3861 2748 3925 2752
rect 3861 2692 3865 2748
rect 3865 2692 3921 2748
rect 3921 2692 3925 2748
rect 3861 2688 3925 2692
rect 3941 2748 4005 2752
rect 3941 2692 3945 2748
rect 3945 2692 4001 2748
rect 4001 2692 4005 2748
rect 3941 2688 4005 2692
rect 4021 2748 4085 2752
rect 4021 2692 4025 2748
rect 4025 2692 4081 2748
rect 4081 2692 4085 2748
rect 4021 2688 4085 2692
rect 5667 2748 5731 2752
rect 5667 2692 5671 2748
rect 5671 2692 5727 2748
rect 5727 2692 5731 2748
rect 5667 2688 5731 2692
rect 5747 2748 5811 2752
rect 5747 2692 5751 2748
rect 5751 2692 5807 2748
rect 5807 2692 5811 2748
rect 5747 2688 5811 2692
rect 5827 2748 5891 2752
rect 5827 2692 5831 2748
rect 5831 2692 5887 2748
rect 5887 2692 5891 2748
rect 5827 2688 5891 2692
rect 5907 2748 5971 2752
rect 5907 2692 5911 2748
rect 5911 2692 5967 2748
rect 5967 2692 5971 2748
rect 5907 2688 5971 2692
rect 7553 2748 7617 2752
rect 7553 2692 7557 2748
rect 7557 2692 7613 2748
rect 7613 2692 7617 2748
rect 7553 2688 7617 2692
rect 7633 2748 7697 2752
rect 7633 2692 7637 2748
rect 7637 2692 7693 2748
rect 7693 2692 7697 2748
rect 7633 2688 7697 2692
rect 7713 2748 7777 2752
rect 7713 2692 7717 2748
rect 7717 2692 7773 2748
rect 7773 2692 7777 2748
rect 7713 2688 7777 2692
rect 7793 2748 7857 2752
rect 7793 2692 7797 2748
rect 7797 2692 7853 2748
rect 7853 2692 7857 2748
rect 7793 2688 7857 2692
rect 2555 2204 2619 2208
rect 2555 2148 2559 2204
rect 2559 2148 2615 2204
rect 2615 2148 2619 2204
rect 2555 2144 2619 2148
rect 2635 2204 2699 2208
rect 2635 2148 2639 2204
rect 2639 2148 2695 2204
rect 2695 2148 2699 2204
rect 2635 2144 2699 2148
rect 2715 2204 2779 2208
rect 2715 2148 2719 2204
rect 2719 2148 2775 2204
rect 2775 2148 2779 2204
rect 2715 2144 2779 2148
rect 2795 2204 2859 2208
rect 2795 2148 2799 2204
rect 2799 2148 2855 2204
rect 2855 2148 2859 2204
rect 2795 2144 2859 2148
rect 4441 2204 4505 2208
rect 4441 2148 4445 2204
rect 4445 2148 4501 2204
rect 4501 2148 4505 2204
rect 4441 2144 4505 2148
rect 4521 2204 4585 2208
rect 4521 2148 4525 2204
rect 4525 2148 4581 2204
rect 4581 2148 4585 2204
rect 4521 2144 4585 2148
rect 4601 2204 4665 2208
rect 4601 2148 4605 2204
rect 4605 2148 4661 2204
rect 4661 2148 4665 2204
rect 4601 2144 4665 2148
rect 4681 2204 4745 2208
rect 4681 2148 4685 2204
rect 4685 2148 4741 2204
rect 4741 2148 4745 2204
rect 4681 2144 4745 2148
rect 6327 2204 6391 2208
rect 6327 2148 6331 2204
rect 6331 2148 6387 2204
rect 6387 2148 6391 2204
rect 6327 2144 6391 2148
rect 6407 2204 6471 2208
rect 6407 2148 6411 2204
rect 6411 2148 6467 2204
rect 6467 2148 6471 2204
rect 6407 2144 6471 2148
rect 6487 2204 6551 2208
rect 6487 2148 6491 2204
rect 6491 2148 6547 2204
rect 6547 2148 6551 2204
rect 6487 2144 6551 2148
rect 6567 2204 6631 2208
rect 6567 2148 6571 2204
rect 6571 2148 6627 2204
rect 6627 2148 6631 2204
rect 6567 2144 6631 2148
rect 8213 2204 8277 2208
rect 8213 2148 8217 2204
rect 8217 2148 8273 2204
rect 8273 2148 8277 2204
rect 8213 2144 8277 2148
rect 8293 2204 8357 2208
rect 8293 2148 8297 2204
rect 8297 2148 8353 2204
rect 8353 2148 8357 2204
rect 8293 2144 8357 2148
rect 8373 2204 8437 2208
rect 8373 2148 8377 2204
rect 8377 2148 8433 2204
rect 8433 2148 8437 2204
rect 8373 2144 8437 2148
rect 8453 2204 8517 2208
rect 8453 2148 8457 2204
rect 8457 2148 8513 2204
rect 8513 2148 8517 2204
rect 8453 2144 8517 2148
<< metal4 >>
rect 1887 9280 2207 9296
rect 1887 9216 1895 9280
rect 1959 9216 1975 9280
rect 2039 9216 2055 9280
rect 2119 9216 2135 9280
rect 2199 9216 2207 9280
rect 1887 8482 2207 9216
rect 1887 8246 1929 8482
rect 2165 8246 2207 8482
rect 1887 8192 2207 8246
rect 1887 8128 1895 8192
rect 1959 8128 1975 8192
rect 2039 8128 2055 8192
rect 2119 8128 2135 8192
rect 2199 8128 2207 8192
rect 1887 7104 2207 8128
rect 1887 7040 1895 7104
rect 1959 7040 1975 7104
rect 2039 7040 2055 7104
rect 2119 7040 2135 7104
rect 2199 7040 2207 7104
rect 1887 6714 2207 7040
rect 1887 6478 1929 6714
rect 2165 6478 2207 6714
rect 1887 6016 2207 6478
rect 1887 5952 1895 6016
rect 1959 5952 1975 6016
rect 2039 5952 2055 6016
rect 2119 5952 2135 6016
rect 2199 5952 2207 6016
rect 1887 4946 2207 5952
rect 1887 4928 1929 4946
rect 2165 4928 2207 4946
rect 1887 4864 1895 4928
rect 2199 4864 2207 4928
rect 1887 4710 1929 4864
rect 2165 4710 2207 4864
rect 1887 3840 2207 4710
rect 1887 3776 1895 3840
rect 1959 3776 1975 3840
rect 2039 3776 2055 3840
rect 2119 3776 2135 3840
rect 2199 3776 2207 3840
rect 1887 3178 2207 3776
rect 1887 2942 1929 3178
rect 2165 2942 2207 3178
rect 1887 2752 2207 2942
rect 1887 2688 1895 2752
rect 1959 2688 1975 2752
rect 2039 2688 2055 2752
rect 2119 2688 2135 2752
rect 2199 2688 2207 2752
rect 1887 2128 2207 2688
rect 2547 9142 2867 9296
rect 2547 8906 2589 9142
rect 2825 8906 2867 9142
rect 2547 8736 2867 8906
rect 2547 8672 2555 8736
rect 2619 8672 2635 8736
rect 2699 8672 2715 8736
rect 2779 8672 2795 8736
rect 2859 8672 2867 8736
rect 2547 7648 2867 8672
rect 2547 7584 2555 7648
rect 2619 7584 2635 7648
rect 2699 7584 2715 7648
rect 2779 7584 2795 7648
rect 2859 7584 2867 7648
rect 2547 7374 2867 7584
rect 2547 7138 2589 7374
rect 2825 7138 2867 7374
rect 2547 6560 2867 7138
rect 2547 6496 2555 6560
rect 2619 6496 2635 6560
rect 2699 6496 2715 6560
rect 2779 6496 2795 6560
rect 2859 6496 2867 6560
rect 2547 5606 2867 6496
rect 2547 5472 2589 5606
rect 2825 5472 2867 5606
rect 2547 5408 2555 5472
rect 2859 5408 2867 5472
rect 2547 5370 2589 5408
rect 2825 5370 2867 5408
rect 2547 4384 2867 5370
rect 2547 4320 2555 4384
rect 2619 4320 2635 4384
rect 2699 4320 2715 4384
rect 2779 4320 2795 4384
rect 2859 4320 2867 4384
rect 2547 3838 2867 4320
rect 2547 3602 2589 3838
rect 2825 3602 2867 3838
rect 2547 3296 2867 3602
rect 2547 3232 2555 3296
rect 2619 3232 2635 3296
rect 2699 3232 2715 3296
rect 2779 3232 2795 3296
rect 2859 3232 2867 3296
rect 2547 2208 2867 3232
rect 2547 2144 2555 2208
rect 2619 2144 2635 2208
rect 2699 2144 2715 2208
rect 2779 2144 2795 2208
rect 2859 2144 2867 2208
rect 2547 2128 2867 2144
rect 3773 9280 4093 9296
rect 3773 9216 3781 9280
rect 3845 9216 3861 9280
rect 3925 9216 3941 9280
rect 4005 9216 4021 9280
rect 4085 9216 4093 9280
rect 3773 8482 4093 9216
rect 3773 8246 3815 8482
rect 4051 8246 4093 8482
rect 3773 8192 4093 8246
rect 3773 8128 3781 8192
rect 3845 8128 3861 8192
rect 3925 8128 3941 8192
rect 4005 8128 4021 8192
rect 4085 8128 4093 8192
rect 3773 7104 4093 8128
rect 3773 7040 3781 7104
rect 3845 7040 3861 7104
rect 3925 7040 3941 7104
rect 4005 7040 4021 7104
rect 4085 7040 4093 7104
rect 3773 6714 4093 7040
rect 3773 6478 3815 6714
rect 4051 6478 4093 6714
rect 3773 6016 4093 6478
rect 3773 5952 3781 6016
rect 3845 5952 3861 6016
rect 3925 5952 3941 6016
rect 4005 5952 4021 6016
rect 4085 5952 4093 6016
rect 3773 4946 4093 5952
rect 3773 4928 3815 4946
rect 4051 4928 4093 4946
rect 3773 4864 3781 4928
rect 4085 4864 4093 4928
rect 3773 4710 3815 4864
rect 4051 4710 4093 4864
rect 3773 3840 4093 4710
rect 3773 3776 3781 3840
rect 3845 3776 3861 3840
rect 3925 3776 3941 3840
rect 4005 3776 4021 3840
rect 4085 3776 4093 3840
rect 3773 3178 4093 3776
rect 3773 2942 3815 3178
rect 4051 2942 4093 3178
rect 3773 2752 4093 2942
rect 3773 2688 3781 2752
rect 3845 2688 3861 2752
rect 3925 2688 3941 2752
rect 4005 2688 4021 2752
rect 4085 2688 4093 2752
rect 3773 2128 4093 2688
rect 4433 9142 4753 9296
rect 4433 8906 4475 9142
rect 4711 8906 4753 9142
rect 4433 8736 4753 8906
rect 4433 8672 4441 8736
rect 4505 8672 4521 8736
rect 4585 8672 4601 8736
rect 4665 8672 4681 8736
rect 4745 8672 4753 8736
rect 4433 7648 4753 8672
rect 4433 7584 4441 7648
rect 4505 7584 4521 7648
rect 4585 7584 4601 7648
rect 4665 7584 4681 7648
rect 4745 7584 4753 7648
rect 4433 7374 4753 7584
rect 4433 7138 4475 7374
rect 4711 7138 4753 7374
rect 4433 6560 4753 7138
rect 4433 6496 4441 6560
rect 4505 6496 4521 6560
rect 4585 6496 4601 6560
rect 4665 6496 4681 6560
rect 4745 6496 4753 6560
rect 4433 5606 4753 6496
rect 4433 5472 4475 5606
rect 4711 5472 4753 5606
rect 4433 5408 4441 5472
rect 4745 5408 4753 5472
rect 4433 5370 4475 5408
rect 4711 5370 4753 5408
rect 4433 4384 4753 5370
rect 4433 4320 4441 4384
rect 4505 4320 4521 4384
rect 4585 4320 4601 4384
rect 4665 4320 4681 4384
rect 4745 4320 4753 4384
rect 4433 3838 4753 4320
rect 4433 3602 4475 3838
rect 4711 3602 4753 3838
rect 4433 3296 4753 3602
rect 4433 3232 4441 3296
rect 4505 3232 4521 3296
rect 4585 3232 4601 3296
rect 4665 3232 4681 3296
rect 4745 3232 4753 3296
rect 4433 2208 4753 3232
rect 4433 2144 4441 2208
rect 4505 2144 4521 2208
rect 4585 2144 4601 2208
rect 4665 2144 4681 2208
rect 4745 2144 4753 2208
rect 4433 2128 4753 2144
rect 5659 9280 5979 9296
rect 5659 9216 5667 9280
rect 5731 9216 5747 9280
rect 5811 9216 5827 9280
rect 5891 9216 5907 9280
rect 5971 9216 5979 9280
rect 5659 8482 5979 9216
rect 5659 8246 5701 8482
rect 5937 8246 5979 8482
rect 5659 8192 5979 8246
rect 5659 8128 5667 8192
rect 5731 8128 5747 8192
rect 5811 8128 5827 8192
rect 5891 8128 5907 8192
rect 5971 8128 5979 8192
rect 5659 7104 5979 8128
rect 5659 7040 5667 7104
rect 5731 7040 5747 7104
rect 5811 7040 5827 7104
rect 5891 7040 5907 7104
rect 5971 7040 5979 7104
rect 5659 6714 5979 7040
rect 5659 6478 5701 6714
rect 5937 6478 5979 6714
rect 5659 6016 5979 6478
rect 5659 5952 5667 6016
rect 5731 5952 5747 6016
rect 5811 5952 5827 6016
rect 5891 5952 5907 6016
rect 5971 5952 5979 6016
rect 5659 4946 5979 5952
rect 5659 4928 5701 4946
rect 5937 4928 5979 4946
rect 5659 4864 5667 4928
rect 5971 4864 5979 4928
rect 5659 4710 5701 4864
rect 5937 4710 5979 4864
rect 5659 3840 5979 4710
rect 5659 3776 5667 3840
rect 5731 3776 5747 3840
rect 5811 3776 5827 3840
rect 5891 3776 5907 3840
rect 5971 3776 5979 3840
rect 5659 3178 5979 3776
rect 5659 2942 5701 3178
rect 5937 2942 5979 3178
rect 5659 2752 5979 2942
rect 5659 2688 5667 2752
rect 5731 2688 5747 2752
rect 5811 2688 5827 2752
rect 5891 2688 5907 2752
rect 5971 2688 5979 2752
rect 5659 2128 5979 2688
rect 6319 9142 6639 9296
rect 6319 8906 6361 9142
rect 6597 8906 6639 9142
rect 6319 8736 6639 8906
rect 6319 8672 6327 8736
rect 6391 8672 6407 8736
rect 6471 8672 6487 8736
rect 6551 8672 6567 8736
rect 6631 8672 6639 8736
rect 6319 7648 6639 8672
rect 6319 7584 6327 7648
rect 6391 7584 6407 7648
rect 6471 7584 6487 7648
rect 6551 7584 6567 7648
rect 6631 7584 6639 7648
rect 6319 7374 6639 7584
rect 6319 7138 6361 7374
rect 6597 7138 6639 7374
rect 6319 6560 6639 7138
rect 6319 6496 6327 6560
rect 6391 6496 6407 6560
rect 6471 6496 6487 6560
rect 6551 6496 6567 6560
rect 6631 6496 6639 6560
rect 6319 5606 6639 6496
rect 6319 5472 6361 5606
rect 6597 5472 6639 5606
rect 6319 5408 6327 5472
rect 6631 5408 6639 5472
rect 6319 5370 6361 5408
rect 6597 5370 6639 5408
rect 6319 4384 6639 5370
rect 6319 4320 6327 4384
rect 6391 4320 6407 4384
rect 6471 4320 6487 4384
rect 6551 4320 6567 4384
rect 6631 4320 6639 4384
rect 6319 3838 6639 4320
rect 6319 3602 6361 3838
rect 6597 3602 6639 3838
rect 6319 3296 6639 3602
rect 6319 3232 6327 3296
rect 6391 3232 6407 3296
rect 6471 3232 6487 3296
rect 6551 3232 6567 3296
rect 6631 3232 6639 3296
rect 6319 2208 6639 3232
rect 6319 2144 6327 2208
rect 6391 2144 6407 2208
rect 6471 2144 6487 2208
rect 6551 2144 6567 2208
rect 6631 2144 6639 2208
rect 6319 2128 6639 2144
rect 7545 9280 7865 9296
rect 7545 9216 7553 9280
rect 7617 9216 7633 9280
rect 7697 9216 7713 9280
rect 7777 9216 7793 9280
rect 7857 9216 7865 9280
rect 7545 8482 7865 9216
rect 7545 8246 7587 8482
rect 7823 8246 7865 8482
rect 7545 8192 7865 8246
rect 7545 8128 7553 8192
rect 7617 8128 7633 8192
rect 7697 8128 7713 8192
rect 7777 8128 7793 8192
rect 7857 8128 7865 8192
rect 7545 7104 7865 8128
rect 7545 7040 7553 7104
rect 7617 7040 7633 7104
rect 7697 7040 7713 7104
rect 7777 7040 7793 7104
rect 7857 7040 7865 7104
rect 7545 6714 7865 7040
rect 7545 6478 7587 6714
rect 7823 6478 7865 6714
rect 7545 6016 7865 6478
rect 7545 5952 7553 6016
rect 7617 5952 7633 6016
rect 7697 5952 7713 6016
rect 7777 5952 7793 6016
rect 7857 5952 7865 6016
rect 7545 4946 7865 5952
rect 7545 4928 7587 4946
rect 7823 4928 7865 4946
rect 7545 4864 7553 4928
rect 7857 4864 7865 4928
rect 7545 4710 7587 4864
rect 7823 4710 7865 4864
rect 7545 3840 7865 4710
rect 7545 3776 7553 3840
rect 7617 3776 7633 3840
rect 7697 3776 7713 3840
rect 7777 3776 7793 3840
rect 7857 3776 7865 3840
rect 7545 3178 7865 3776
rect 7545 2942 7587 3178
rect 7823 2942 7865 3178
rect 7545 2752 7865 2942
rect 7545 2688 7553 2752
rect 7617 2688 7633 2752
rect 7697 2688 7713 2752
rect 7777 2688 7793 2752
rect 7857 2688 7865 2752
rect 7545 2128 7865 2688
rect 8205 9142 8525 9296
rect 8205 8906 8247 9142
rect 8483 8906 8525 9142
rect 8205 8736 8525 8906
rect 8205 8672 8213 8736
rect 8277 8672 8293 8736
rect 8357 8672 8373 8736
rect 8437 8672 8453 8736
rect 8517 8672 8525 8736
rect 8205 7648 8525 8672
rect 8205 7584 8213 7648
rect 8277 7584 8293 7648
rect 8357 7584 8373 7648
rect 8437 7584 8453 7648
rect 8517 7584 8525 7648
rect 8205 7374 8525 7584
rect 8205 7138 8247 7374
rect 8483 7138 8525 7374
rect 8205 6560 8525 7138
rect 8205 6496 8213 6560
rect 8277 6496 8293 6560
rect 8357 6496 8373 6560
rect 8437 6496 8453 6560
rect 8517 6496 8525 6560
rect 8205 5606 8525 6496
rect 8205 5472 8247 5606
rect 8483 5472 8525 5606
rect 8205 5408 8213 5472
rect 8517 5408 8525 5472
rect 8205 5370 8247 5408
rect 8483 5370 8525 5408
rect 8205 4384 8525 5370
rect 8205 4320 8213 4384
rect 8277 4320 8293 4384
rect 8357 4320 8373 4384
rect 8437 4320 8453 4384
rect 8517 4320 8525 4384
rect 8205 3838 8525 4320
rect 8205 3602 8247 3838
rect 8483 3602 8525 3838
rect 8205 3296 8525 3602
rect 8205 3232 8213 3296
rect 8277 3232 8293 3296
rect 8357 3232 8373 3296
rect 8437 3232 8453 3296
rect 8517 3232 8525 3296
rect 8205 2208 8525 3232
rect 8205 2144 8213 2208
rect 8277 2144 8293 2208
rect 8357 2144 8373 2208
rect 8437 2144 8453 2208
rect 8517 2144 8525 2208
rect 8205 2128 8525 2144
<< via4 >>
rect 1929 8246 2165 8482
rect 1929 6478 2165 6714
rect 1929 4928 2165 4946
rect 1929 4864 1959 4928
rect 1959 4864 1975 4928
rect 1975 4864 2039 4928
rect 2039 4864 2055 4928
rect 2055 4864 2119 4928
rect 2119 4864 2135 4928
rect 2135 4864 2165 4928
rect 1929 4710 2165 4864
rect 1929 2942 2165 3178
rect 2589 8906 2825 9142
rect 2589 7138 2825 7374
rect 2589 5472 2825 5606
rect 2589 5408 2619 5472
rect 2619 5408 2635 5472
rect 2635 5408 2699 5472
rect 2699 5408 2715 5472
rect 2715 5408 2779 5472
rect 2779 5408 2795 5472
rect 2795 5408 2825 5472
rect 2589 5370 2825 5408
rect 2589 3602 2825 3838
rect 3815 8246 4051 8482
rect 3815 6478 4051 6714
rect 3815 4928 4051 4946
rect 3815 4864 3845 4928
rect 3845 4864 3861 4928
rect 3861 4864 3925 4928
rect 3925 4864 3941 4928
rect 3941 4864 4005 4928
rect 4005 4864 4021 4928
rect 4021 4864 4051 4928
rect 3815 4710 4051 4864
rect 3815 2942 4051 3178
rect 4475 8906 4711 9142
rect 4475 7138 4711 7374
rect 4475 5472 4711 5606
rect 4475 5408 4505 5472
rect 4505 5408 4521 5472
rect 4521 5408 4585 5472
rect 4585 5408 4601 5472
rect 4601 5408 4665 5472
rect 4665 5408 4681 5472
rect 4681 5408 4711 5472
rect 4475 5370 4711 5408
rect 4475 3602 4711 3838
rect 5701 8246 5937 8482
rect 5701 6478 5937 6714
rect 5701 4928 5937 4946
rect 5701 4864 5731 4928
rect 5731 4864 5747 4928
rect 5747 4864 5811 4928
rect 5811 4864 5827 4928
rect 5827 4864 5891 4928
rect 5891 4864 5907 4928
rect 5907 4864 5937 4928
rect 5701 4710 5937 4864
rect 5701 2942 5937 3178
rect 6361 8906 6597 9142
rect 6361 7138 6597 7374
rect 6361 5472 6597 5606
rect 6361 5408 6391 5472
rect 6391 5408 6407 5472
rect 6407 5408 6471 5472
rect 6471 5408 6487 5472
rect 6487 5408 6551 5472
rect 6551 5408 6567 5472
rect 6567 5408 6597 5472
rect 6361 5370 6597 5408
rect 6361 3602 6597 3838
rect 7587 8246 7823 8482
rect 7587 6478 7823 6714
rect 7587 4928 7823 4946
rect 7587 4864 7617 4928
rect 7617 4864 7633 4928
rect 7633 4864 7697 4928
rect 7697 4864 7713 4928
rect 7713 4864 7777 4928
rect 7777 4864 7793 4928
rect 7793 4864 7823 4928
rect 7587 4710 7823 4864
rect 7587 2942 7823 3178
rect 8247 8906 8483 9142
rect 8247 7138 8483 7374
rect 8247 5472 8483 5606
rect 8247 5408 8277 5472
rect 8277 5408 8293 5472
rect 8293 5408 8357 5472
rect 8357 5408 8373 5472
rect 8373 5408 8437 5472
rect 8437 5408 8453 5472
rect 8453 5408 8483 5472
rect 8247 5370 8483 5408
rect 8247 3602 8483 3838
<< metal5 >>
rect 1056 9142 8696 9184
rect 1056 8906 2589 9142
rect 2825 8906 4475 9142
rect 4711 8906 6361 9142
rect 6597 8906 8247 9142
rect 8483 8906 8696 9142
rect 1056 8864 8696 8906
rect 1056 8482 8696 8524
rect 1056 8246 1929 8482
rect 2165 8246 3815 8482
rect 4051 8246 5701 8482
rect 5937 8246 7587 8482
rect 7823 8246 8696 8482
rect 1056 8204 8696 8246
rect 1056 7374 8696 7416
rect 1056 7138 2589 7374
rect 2825 7138 4475 7374
rect 4711 7138 6361 7374
rect 6597 7138 8247 7374
rect 8483 7138 8696 7374
rect 1056 7096 8696 7138
rect 1056 6714 8696 6756
rect 1056 6478 1929 6714
rect 2165 6478 3815 6714
rect 4051 6478 5701 6714
rect 5937 6478 7587 6714
rect 7823 6478 8696 6714
rect 1056 6436 8696 6478
rect 1056 5606 8696 5648
rect 1056 5370 2589 5606
rect 2825 5370 4475 5606
rect 4711 5370 6361 5606
rect 6597 5370 8247 5606
rect 8483 5370 8696 5606
rect 1056 5328 8696 5370
rect 1056 4946 8696 4988
rect 1056 4710 1929 4946
rect 2165 4710 3815 4946
rect 4051 4710 5701 4946
rect 5937 4710 7587 4946
rect 7823 4710 8696 4946
rect 1056 4668 8696 4710
rect 1056 3838 8696 3880
rect 1056 3602 2589 3838
rect 2825 3602 4475 3838
rect 4711 3602 6361 3838
rect 6597 3602 8247 3838
rect 8483 3602 8696 3838
rect 1056 3560 8696 3602
rect 1056 3178 8696 3220
rect 1056 2942 1929 3178
rect 2165 2942 3815 3178
rect 4051 2942 5701 3178
rect 5937 2942 7587 3178
rect 7823 2942 8696 3178
rect 1056 2900 8696 2942
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1670211287
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35
timestamp 1670211287
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1670211287
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1670211287
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1670211287
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1670211287
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1670211287
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1670211287
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1670211287
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1670211287
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1670211287
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1670211287
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1670211287
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1670211287
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1670211287
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1670211287
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1670211287
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1670211287
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1670211287
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1670211287
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1670211287
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1670211287
transform 1 0 8188 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1670211287
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1670211287
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1670211287
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_36
timestamp 1670211287
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1670211287
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1670211287
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1670211287
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1670211287
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1670211287
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1670211287
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1670211287
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1670211287
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_29
timestamp 1670211287
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_35
timestamp 1670211287
transform 1 0 4324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1670211287
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_60
timestamp 1670211287
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_72
timestamp 1670211287
transform 1 0 7728 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_78
timestamp 1670211287
transform 1 0 8280 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1670211287
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1670211287
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1670211287
transform 1 0 2852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_25
timestamp 1670211287
transform 1 0 3404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1670211287
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_46
timestamp 1670211287
transform 1 0 5336 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1670211287
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1670211287
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_75
timestamp 1670211287
transform 1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1670211287
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_15
timestamp 1670211287
transform 1 0 2484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_21
timestamp 1670211287
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1670211287
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_37
timestamp 1670211287
transform 1 0 4508 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1670211287
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_54
timestamp 1670211287
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_66
timestamp 1670211287
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_78
timestamp 1670211287
transform 1 0 8280 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1670211287
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1670211287
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1670211287
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 1670211287
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_38
timestamp 1670211287
transform 1 0 4600 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1670211287
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1670211287
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_62
timestamp 1670211287
transform 1 0 6808 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1670211287
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1670211287
transform 1 0 8280 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1670211287
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_8
timestamp 1670211287
transform 1 0 1840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1670211287
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1670211287
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_39
timestamp 1670211287
transform 1 0 4692 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_63
timestamp 1670211287
transform 1 0 6900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_75
timestamp 1670211287
transform 1 0 8004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1670211287
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1670211287
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1670211287
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1670211287
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1670211287
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_75
timestamp 1670211287
transform 1 0 8004 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1670211287
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1670211287
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1670211287
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1670211287
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1670211287
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_37
timestamp 1670211287
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_44
timestamp 1670211287
transform 1 0 5152 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_56
timestamp 1670211287
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1670211287
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_72
timestamp 1670211287
transform 1 0 7728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 1670211287
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1670211287
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_9
timestamp 1670211287
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_21
timestamp 1670211287
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_33
timestamp 1670211287
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp 1670211287
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1670211287
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1670211287
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_69
timestamp 1670211287
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1670211287
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1670211287
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1670211287
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1670211287
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1670211287
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1670211287
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1670211287
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_53
timestamp 1670211287
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1670211287
transform 1 0 6348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_63
timestamp 1670211287
transform 1 0 6900 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp 1670211287
transform 1 0 7636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1670211287
transform 1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1670211287
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1670211287
transform -1 0 8648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1670211287
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1670211287
transform -1 0 8648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1670211287
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1670211287
transform -1 0 8648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1670211287
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1670211287
transform -1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1670211287
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1670211287
transform -1 0 8648 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1670211287
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1670211287
transform -1 0 8648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1670211287
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1670211287
transform -1 0 8648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1670211287
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1670211287
transform -1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1670211287
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1670211287
transform -1 0 8648 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1670211287
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1670211287
transform -1 0 8648 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1670211287
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1670211287
transform -1 0 8648 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1670211287
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1670211287
transform -1 0 8648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1670211287
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1670211287
transform -1 0 8648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1670211287
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1670211287
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1670211287
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1670211287
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1670211287
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1670211287
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1670211287
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1670211287
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1670211287
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1670211287
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1670211287
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1670211287
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1670211287
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1670211287
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 3128 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform -1 0 3404 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform -1 0 4416 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 4048 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 3956 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform -1 0 3496 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _25_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 4876 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform -1 0 6072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform -1 0 5888 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _28_
timestamp 1670211287
transform -1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _29_
timestamp 1670211287
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _30_
timestamp 1670211287
transform 1 0 4784 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _31_
timestamp 1670211287
transform -1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 4048 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1670211287
transform 1 0 4232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _34_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 6532 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _35_
timestamp 1670211287
transform 1 0 2944 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _36_
timestamp 1670211287
transform -1 0 3036 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _37_
timestamp 1670211287
transform 1 0 5428 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _38_
timestamp 1670211287
transform 1 0 6532 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 4416 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _40_
timestamp 1670211287
transform 1 0 4140 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1670211287
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1670211287
transform -1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670211287
transform 1 0 7820 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1670211287
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1670211287
transform 1 0 6532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1670211287
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1670211287
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1670211287
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1670211287
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1670211287
transform 1 0 1564 0 1 8704
box -38 -48 406 592
<< labels >>
flabel metal4 s 2547 2128 2867 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4433 2128 4753 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6319 2128 6639 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8205 2128 8525 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3560 8696 3880 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5328 8696 5648 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7096 8696 7416 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8864 8696 9184 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1887 2128 2207 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3773 2128 4093 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5659 2128 5979 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7545 2128 7865 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 2900 8696 3220 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4668 8696 4988 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 6436 8696 6756 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8204 8696 8524 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9678 11122 9734 11922 0 FreeSans 224 90 0 0 bcd_value[0]
port 2 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 bcd_value[1]
port 3 nsew signal tristate
flabel metal2 s 5814 11122 5870 11922 0 FreeSans 224 90 0 0 bcd_value[2]
port 4 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 bcd_value[3]
port 5 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 clk
port 6 nsew signal input
flabel metal3 s 8978 7488 9778 7608 0 FreeSans 480 0 0 0 gray_count[0]
port 7 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gray_count[1]
port 8 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 gray_count[2]
port 9 nsew signal tristate
flabel metal2 s 1306 11122 1362 11922 0 FreeSans 224 90 0 0 gray_count[3]
port 10 nsew signal tristate
flabel metal3 s 8978 2728 9778 2848 0 FreeSans 480 0 0 0 rst
port 11 nsew signal input
rlabel metal1 4876 8704 4876 8704 0 VGND
rlabel metal1 4876 9248 4876 9248 0 VPWR
rlabel metal1 6762 6426 6762 6426 0 _00_
rlabel via1 3261 4182 3261 4182 0 _01_
rlabel metal1 3000 7378 3000 7378 0 _02_
rlabel metal2 5842 6562 5842 6562 0 _03_
rlabel metal1 6624 4794 6624 4794 0 _04_
rlabel via1 4733 4590 4733 4590 0 _05_
rlabel metal1 4354 7446 4354 7446 0 _06_
rlabel metal2 4002 5270 4002 5270 0 _07_
rlabel metal1 3496 5338 3496 5338 0 _08_
rlabel metal2 3450 4794 3450 4794 0 _09_
rlabel metal1 4462 6800 4462 6800 0 _10_
rlabel metal1 3726 6766 3726 6766 0 _11_
rlabel via1 5290 6290 5290 6290 0 _12_
rlabel metal1 5842 6290 5842 6290 0 _13_
rlabel metal1 5106 5202 5106 5202 0 _14_
rlabel metal1 4646 5678 4646 5678 0 _15_
rlabel metal1 4416 5882 4416 5882 0 _16_
rlabel metal1 8740 9146 8740 9146 0 bcd_value[0]
rlabel metal2 46 1520 46 1520 0 bcd_value[1]
rlabel metal1 6486 9146 6486 9146 0 bcd_value[2]
rlabel metal2 8418 1095 8418 1095 0 bcd_value[3]
rlabel metal3 1188 4148 1188 4148 0 clk
rlabel metal2 8050 7565 8050 7565 0 gray_count[0]
rlabel metal2 3910 1520 3910 1520 0 gray_count[1]
rlabel metal2 1794 8755 1794 8755 0 gray_count[2]
rlabel metal1 1564 9146 1564 9146 0 gray_count[3]
rlabel metal2 2990 4318 2990 4318 0 net1
rlabel metal1 1564 6630 1564 6630 0 net10
rlabel metal1 6670 4590 6670 4590 0 net2
rlabel metal2 3174 5440 3174 5440 0 net3
rlabel metal2 3174 3706 3174 3706 0 net4
rlabel metal1 5352 5610 5352 5610 0 net5
rlabel metal1 2438 6698 2438 6698 0 net6
rlabel metal2 7958 7684 7958 7684 0 net7
rlabel metal2 4278 3162 4278 3162 0 net8
rlabel metal2 1610 7990 1610 7990 0 net9
rlabel metal2 8050 2907 8050 2907 0 rst
<< properties >>
string FIXED_BBOX 0 0 9778 11922
<< end >>

* NGSPICE file created from iiitb_gray_cntr.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

.subckt iiitb_gray_cntr VGND VPWR bcd_value[0] bcd_value[1] bcd_value[2] bcd_value[3]
+ clk gray_count[0] gray_count[1] gray_count[2] gray_count[3] rst
XFILLER_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput7 net7 VGND VGND VPWR VPWR gray_count[0] sky130_fd_sc_hd__buf_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput10 net10 VGND VGND VPWR VPWR gray_count[3] sky130_fd_sc_hd__buf_2
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput8 net8 VGND VGND VPWR VPWR gray_count[1] sky130_fd_sc_hd__buf_2
XFILLER_3_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR gray_count[2] sky130_fd_sc_hd__buf_2
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29_ net3 net4 net2 VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28_ net3 net2 VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__nor2_1
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27_ net6 _12_ _13_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__o21a_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26_ net6 _12_ net2 VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25_ net3 net4 net5 VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__and3_1
XFILLER_7_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24_ net6 _10_ _11_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__a21boi_1
X_41_ net6 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_40_ net1 _06_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23_ net6 _10_ net2 VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__o21ba_1
XFILLER_11_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22_ net3 net4 net5 VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__a21o_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21_ _09_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__clkbuf_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 clk VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_20_ net2 _07_ _08_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__and3b_1
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 rst VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_39_ net1 _05_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfxtp_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_38_ net1 _04_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_37_ net1 _03_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36_ net1 _02_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfxtp_1
X_19_ net3 net4 net5 VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__or3_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35_ net1 _01_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfxtp_1
X_18_ net3 net4 net5 VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__o21ai_1
XTAP_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34_ net1 _00_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfxtp_1
X_17_ net4 net2 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33_ _16_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ _10_ _15_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__and2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31_ net2 _12_ VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__nor2_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30_ net3 net4 _14_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__o21a_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput3 net3 VGND VGND VPWR VPWR bcd_value[0] sky130_fd_sc_hd__buf_2
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput4 net4 VGND VGND VPWR VPWR bcd_value[1] sky130_fd_sc_hd__buf_2
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput5 net5 VGND VGND VPWR VPWR bcd_value[2] sky130_fd_sc_hd__buf_2
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput6 net6 VGND VGND VPWR VPWR bcd_value[3] sky130_fd_sc_hd__buf_2
.ends


magic
tech sky130A
magscale 1 2
timestamp 1670837675
<< obsli1 >>
rect 1104 2159 8648 9265
<< obsm1 >>
rect 14 2128 9462 9296
<< metal2 >>
rect 1306 11122 1362 11922
rect 5814 11122 5870 11922
rect 9678 11122 9734 11922
rect 18 0 74 800
rect 3882 0 3938 800
rect 8390 0 8446 800
<< obsm2 >>
rect 20 11066 1250 11234
rect 1418 11066 5758 11234
rect 5926 11066 9622 11234
rect 20 856 9678 11066
rect 130 800 3826 856
rect 3994 800 8334 856
rect 8502 800 9678 856
<< metal3 >>
rect 0 8848 800 8968
rect 8978 7488 9778 7608
rect 0 4088 800 4208
rect 8978 2728 9778 2848
<< obsm3 >>
rect 800 9048 8978 9281
rect 880 8768 8978 9048
rect 800 7688 8978 8768
rect 800 7408 8898 7688
rect 800 4288 8978 7408
rect 880 4008 8978 4288
rect 800 2928 8978 4008
rect 800 2648 8898 2928
rect 800 2143 8978 2648
<< metal4 >>
rect 1887 2128 2207 9296
rect 2547 2128 2867 9296
rect 3773 2128 4093 9296
rect 4433 2128 4753 9296
rect 5659 2128 5979 9296
rect 6319 2128 6639 9296
rect 7545 2128 7865 9296
rect 8205 2128 8525 9296
<< metal5 >>
rect 1056 8864 8696 9184
rect 1056 8204 8696 8524
rect 1056 7096 8696 7416
rect 1056 6436 8696 6756
rect 1056 5328 8696 5648
rect 1056 4668 8696 4988
rect 1056 3560 8696 3880
rect 1056 2900 8696 3220
<< labels >>
rlabel metal4 s 2547 2128 2867 9296 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4433 2128 4753 9296 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6319 2128 6639 9296 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8205 2128 8525 9296 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3560 8696 3880 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5328 8696 5648 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7096 8696 7416 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8864 8696 9184 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1887 2128 2207 9296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3773 2128 4093 9296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5659 2128 5979 9296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7545 2128 7865 9296 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2900 8696 3220 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4668 8696 4988 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6436 8696 6756 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8204 8696 8524 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 9678 11122 9734 11922 6 bcd_value[0]
port 3 nsew signal output
rlabel metal2 s 18 0 74 800 6 bcd_value[1]
port 4 nsew signal output
rlabel metal2 s 5814 11122 5870 11922 6 bcd_value[2]
port 5 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 bcd_value[3]
port 6 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 clk
port 7 nsew signal input
rlabel metal3 s 8978 7488 9778 7608 6 gray_count[0]
port 8 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 gray_count[1]
port 9 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 gray_count[2]
port 10 nsew signal output
rlabel metal2 s 1306 11122 1362 11922 6 gray_count[3]
port 11 nsew signal output
rlabel metal3 s 8978 2728 9778 2848 6 rst
port 12 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 9778 11922
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 258524
string GDS_FILE /openlane/designs/iiitb_gray_cntr/runs/RUN_2022.12.12_09.32.31/results/signoff/iiitb_gray_cntr.magic.gds
string GDS_START 118870
<< end >>

